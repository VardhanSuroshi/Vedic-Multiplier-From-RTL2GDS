module pes_vedic_mul (a,
    b,
    prod);
 input [7:0] a;
 input [7:0] b;
 output [15:0] prod;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;

 sky130_fd_sc_hd__xor2_1 _314_ (.A(_077_),
    .B(_078_),
    .X(_079_));
 sky130_fd_sc_hd__nor2_1 _315_ (.A(_308_),
    .B(_042_),
    .Y(_080_));
 sky130_fd_sc_hd__nand2_1 _316_ (.A(_011_),
    .B(_080_),
    .Y(_081_));
 sky130_fd_sc_hd__xor2_1 _317_ (.A(_045_),
    .B(_081_),
    .X(_082_));
 sky130_fd_sc_hd__nand2_1 _318_ (.A(_079_),
    .B(_082_),
    .Y(_083_));
 sky130_fd_sc_hd__or2_1 _319_ (.A(_079_),
    .B(_082_),
    .X(_084_));
 sky130_fd_sc_hd__and2_1 _320_ (.A(_083_),
    .B(_084_),
    .X(_085_));
 sky130_fd_sc_hd__o21ai_1 _321_ (.A1(_076_),
    .A2(_049_),
    .B1(_085_),
    .Y(_086_));
 sky130_fd_sc_hd__or3_1 _322_ (.A(_076_),
    .B(_049_),
    .C(_085_),
    .X(_087_));
 sky130_fd_sc_hd__nand2_1 _323_ (.A(_086_),
    .B(_087_),
    .Y(_088_));
 sky130_fd_sc_hd__nand2_1 _324_ (.A(_266_),
    .B(_265_),
    .Y(_089_));
 sky130_fd_sc_hd__or2_1 _325_ (.A(_088_),
    .B(_089_),
    .X(_090_));
 sky130_fd_sc_hd__nand2_1 _326_ (.A(_088_),
    .B(_089_),
    .Y(_091_));
 sky130_fd_sc_hd__nand2_1 _327_ (.A(_090_),
    .B(_091_),
    .Y(_092_));
 sky130_fd_sc_hd__a21oi_1 _328_ (.A1(_053_),
    .A2(_070_),
    .B1(_069_),
    .Y(_093_));
 sky130_fd_sc_hd__or2_1 _329_ (.A(_058_),
    .B(_066_),
    .X(_094_));
 sky130_fd_sc_hd__inv_2 _330_ (.A(_067_),
    .Y(_095_));
 sky130_fd_sc_hd__nand2_1 _331_ (.A(_024_),
    .B(_095_),
    .Y(_096_));
 sky130_fd_sc_hd__buf_2 _332_ (.A(net7),
    .X(_097_));
 sky130_fd_sc_hd__nand2_1 _333_ (.A(_261_),
    .B(_097_),
    .Y(_098_));
 sky130_fd_sc_hd__and3_1 _334_ (.A(_270_),
    .B(_301_),
    .C(_022_),
    .X(_099_));
 sky130_fd_sc_hd__xor2_1 _335_ (.A(_098_),
    .B(_099_),
    .X(_100_));
 sky130_fd_sc_hd__buf_2 _336_ (.A(net8),
    .X(_101_));
 sky130_fd_sc_hd__and3_1 _337_ (.A(_247_),
    .B(_101_),
    .C(_019_),
    .X(_102_));
 sky130_fd_sc_hd__xnor2_1 _338_ (.A(_064_),
    .B(_102_),
    .Y(_103_));
 sky130_fd_sc_hd__nor2_1 _339_ (.A(_100_),
    .B(_103_),
    .Y(_104_));
 sky130_fd_sc_hd__and2_1 _340_ (.A(_100_),
    .B(_103_),
    .X(_105_));
 sky130_fd_sc_hd__or2_1 _341_ (.A(_104_),
    .B(_105_),
    .X(_106_));
 sky130_fd_sc_hd__a21oi_1 _342_ (.A1(_094_),
    .A2(_096_),
    .B1(_106_),
    .Y(_107_));
 sky130_fd_sc_hd__and3_1 _343_ (.A(_094_),
    .B(_096_),
    .C(_106_),
    .X(_108_));
 sky130_fd_sc_hd__nor2_1 _344_ (.A(_107_),
    .B(_108_),
    .Y(_109_));
 sky130_fd_sc_hd__xnor2_1 _345_ (.A(_093_),
    .B(_109_),
    .Y(_110_));
 sky130_fd_sc_hd__xnor2_1 _346_ (.A(_092_),
    .B(_110_),
    .Y(_111_));
 sky130_fd_sc_hd__and2b_1 _347_ (.A_N(_092_),
    .B(_110_),
    .X(_112_));
 sky130_fd_sc_hd__a21o_1 _348_ (.A1(_075_),
    .A2(_111_),
    .B1(_112_),
    .X(_113_));
 sky130_fd_sc_hd__a22o_1 _349_ (.A1(_266_),
    .A2(net14),
    .B1(_265_),
    .B2(_301_),
    .X(_114_));
 sky130_fd_sc_hd__inv_2 _350_ (.A(_301_),
    .Y(_115_));
 sky130_fd_sc_hd__or3_1 _351_ (.A(_115_),
    .B(_042_),
    .C(_089_),
    .X(_116_));
 sky130_fd_sc_hd__nand2_1 _352_ (.A(_114_),
    .B(_116_),
    .Y(_117_));
 sky130_fd_sc_hd__a21o_1 _353_ (.A1(_257_),
    .A2(_265_),
    .B1(_045_),
    .X(_118_));
 sky130_fd_sc_hd__a22o_1 _354_ (.A1(_257_),
    .A2(net16),
    .B1(_038_),
    .B2(_272_),
    .X(_119_));
 sky130_fd_sc_hd__inv_2 _355_ (.A(net16),
    .Y(_120_));
 sky130_fd_sc_hd__or3_1 _356_ (.A(_308_),
    .B(_120_),
    .C(_077_),
    .X(_121_));
 sky130_fd_sc_hd__o2111a_1 _357_ (.A1(_253_),
    .A2(_257_),
    .B1(net16),
    .C1(_038_),
    .D1(_254_),
    .X(_122_));
 sky130_fd_sc_hd__and3_1 _358_ (.A(_119_),
    .B(_121_),
    .C(_122_),
    .X(_123_));
 sky130_fd_sc_hd__a21oi_1 _359_ (.A1(_119_),
    .A2(_121_),
    .B1(_122_),
    .Y(_124_));
 sky130_fd_sc_hd__nor2_1 _360_ (.A(_123_),
    .B(_124_),
    .Y(_125_));
 sky130_fd_sc_hd__a21o_1 _361_ (.A1(_080_),
    .A2(_118_),
    .B1(_125_),
    .X(_126_));
 sky130_fd_sc_hd__nand3_1 _362_ (.A(_080_),
    .B(_125_),
    .C(_118_),
    .Y(_127_));
 sky130_fd_sc_hd__nand2_1 _363_ (.A(_126_),
    .B(_127_),
    .Y(_128_));
 sky130_fd_sc_hd__a21o_1 _364_ (.A1(_084_),
    .A2(_086_),
    .B1(_128_),
    .X(_129_));
 sky130_fd_sc_hd__nand3_1 _365_ (.A(_084_),
    .B(_086_),
    .C(_128_),
    .Y(_130_));
 sky130_fd_sc_hd__and2_1 _366_ (.A(_129_),
    .B(_130_),
    .X(_131_));
 sky130_fd_sc_hd__xor2_1 _367_ (.A(_117_),
    .B(_131_),
    .X(_132_));
 sky130_fd_sc_hd__nor2_1 _368_ (.A(_090_),
    .B(_132_),
    .Y(_133_));
 sky130_fd_sc_hd__and2_1 _369_ (.A(_090_),
    .B(_132_),
    .X(_134_));
 sky130_fd_sc_hd__or2_1 _370_ (.A(_133_),
    .B(_134_),
    .X(_135_));
 sky130_fd_sc_hd__and2b_1 _371_ (.A_N(_093_),
    .B(_109_),
    .X(_136_));
 sky130_fd_sc_hd__a21boi_1 _372_ (.A1(_064_),
    .A2(_102_),
    .B1_N(_062_),
    .Y(_137_));
 sky130_fd_sc_hd__a22o_1 _373_ (.A1(_270_),
    .A2(_097_),
    .B1(_101_),
    .B2(_261_),
    .X(_138_));
 sky130_fd_sc_hd__or3_1 _374_ (.A(_309_),
    .B(_061_),
    .C(_098_),
    .X(_139_));
 sky130_fd_sc_hd__a31o_1 _375_ (.A1(_261_),
    .A2(_097_),
    .A3(_099_),
    .B1(_057_),
    .X(_140_));
 sky130_fd_sc_hd__and3_1 _376_ (.A(_138_),
    .B(_139_),
    .C(_140_),
    .X(_141_));
 sky130_fd_sc_hd__a21oi_1 _377_ (.A1(_138_),
    .A2(_139_),
    .B1(_140_),
    .Y(_142_));
 sky130_fd_sc_hd__or3_1 _378_ (.A(_137_),
    .B(_141_),
    .C(_142_),
    .X(_143_));
 sky130_fd_sc_hd__o21ai_1 _379_ (.A1(_141_),
    .A2(_142_),
    .B1(_137_),
    .Y(_144_));
 sky130_fd_sc_hd__and2_1 _380_ (.A(_143_),
    .B(_144_),
    .X(_145_));
 sky130_fd_sc_hd__o21ai_1 _381_ (.A1(_104_),
    .A2(_107_),
    .B1(_145_),
    .Y(_146_));
 sky130_fd_sc_hd__or3_1 _382_ (.A(_104_),
    .B(_107_),
    .C(_145_),
    .X(_147_));
 sky130_fd_sc_hd__and2_1 _383_ (.A(_146_),
    .B(_147_),
    .X(_148_));
 sky130_fd_sc_hd__xnor2_1 _384_ (.A(_136_),
    .B(_148_),
    .Y(_149_));
 sky130_fd_sc_hd__xor2_1 _385_ (.A(_135_),
    .B(_149_),
    .X(_150_));
 sky130_fd_sc_hd__nor2_1 _386_ (.A(_135_),
    .B(_149_),
    .Y(_151_));
 sky130_fd_sc_hd__a21o_1 _387_ (.A1(_113_),
    .A2(_150_),
    .B1(_151_),
    .X(_152_));
 sky130_fd_sc_hd__and3_1 _388_ (.A(_114_),
    .B(_116_),
    .C(_131_),
    .X(_153_));
 sky130_fd_sc_hd__nand2_1 _389_ (.A(_097_),
    .B(_265_),
    .Y(_154_));
 sky130_fd_sc_hd__and3_1 _390_ (.A(_301_),
    .B(net14),
    .C(_089_),
    .X(_155_));
 sky130_fd_sc_hd__xor2_1 _391_ (.A(_154_),
    .B(_155_),
    .X(_156_));
 sky130_fd_sc_hd__nand2_1 _392_ (.A(_266_),
    .B(_038_),
    .Y(_157_));
 sky130_fd_sc_hd__or2_1 _393_ (.A(_156_),
    .B(_157_),
    .X(_158_));
 sky130_fd_sc_hd__nand2_1 _394_ (.A(_156_),
    .B(_157_),
    .Y(_159_));
 sky130_fd_sc_hd__nand2_1 _395_ (.A(_158_),
    .B(_159_),
    .Y(_160_));
 sky130_fd_sc_hd__a31o_1 _396_ (.A1(_272_),
    .A2(_037_),
    .A3(_077_),
    .B1(_123_),
    .X(_161_));
 sky130_fd_sc_hd__nand3_1 _397_ (.A(_272_),
    .B(_037_),
    .C(_123_),
    .Y(_162_));
 sky130_fd_sc_hd__nand2_1 _398_ (.A(_161_),
    .B(_162_),
    .Y(_163_));
 sky130_fd_sc_hd__a21o_1 _399_ (.A1(_127_),
    .A2(_129_),
    .B1(_163_),
    .X(_164_));
 sky130_fd_sc_hd__nand3_1 _400_ (.A(_127_),
    .B(_129_),
    .C(_163_),
    .Y(_165_));
 sky130_fd_sc_hd__nand2_1 _401_ (.A(_164_),
    .B(_165_),
    .Y(_166_));
 sky130_fd_sc_hd__xor2_1 _402_ (.A(_160_),
    .B(_166_),
    .X(_167_));
 sky130_fd_sc_hd__o21a_1 _403_ (.A1(_153_),
    .A2(_133_),
    .B1(_167_),
    .X(_168_));
 sky130_fd_sc_hd__nor3_1 _404_ (.A(_153_),
    .B(_133_),
    .C(_167_),
    .Y(_169_));
 sky130_fd_sc_hd__nor2_1 _405_ (.A(_168_),
    .B(_169_),
    .Y(_170_));
 sky130_fd_sc_hd__and2_1 _406_ (.A(_136_),
    .B(_148_),
    .X(_171_));
 sky130_fd_sc_hd__and3_1 _407_ (.A(_270_),
    .B(_101_),
    .C(_098_),
    .X(_172_));
 sky130_fd_sc_hd__nor2_1 _408_ (.A(_141_),
    .B(_172_),
    .Y(_173_));
 sky130_fd_sc_hd__a31o_1 _409_ (.A1(_270_),
    .A2(_101_),
    .A3(_141_),
    .B1(_173_),
    .X(_174_));
 sky130_fd_sc_hd__a21o_1 _410_ (.A1(_143_),
    .A2(_146_),
    .B1(_174_),
    .X(_175_));
 sky130_fd_sc_hd__nand3_1 _411_ (.A(_143_),
    .B(_146_),
    .C(_174_),
    .Y(_176_));
 sky130_fd_sc_hd__and2_1 _412_ (.A(_175_),
    .B(_176_),
    .X(_177_));
 sky130_fd_sc_hd__xor2_1 _413_ (.A(_171_),
    .B(_177_),
    .X(_178_));
 sky130_fd_sc_hd__xor2_1 _414_ (.A(_170_),
    .B(_178_),
    .X(_179_));
 sky130_fd_sc_hd__xor2_1 _415_ (.A(_152_),
    .B(_179_),
    .X(net18));
 sky130_fd_sc_hd__and2_1 _416_ (.A(_170_),
    .B(_178_),
    .X(_180_));
 sky130_fd_sc_hd__a21o_1 _417_ (.A1(_152_),
    .A2(_179_),
    .B1(_180_),
    .X(_181_));
 sky130_fd_sc_hd__nor2_1 _418_ (.A(_160_),
    .B(_166_),
    .Y(_182_));
 sky130_fd_sc_hd__a22oi_1 _419_ (.A1(_266_),
    .A2(_037_),
    .B1(_038_),
    .B2(_301_),
    .Y(_183_));
 sky130_fd_sc_hd__and4_1 _420_ (.A(_301_),
    .B(_266_),
    .C(_037_),
    .D(_038_),
    .X(_184_));
 sky130_fd_sc_hd__or2_1 _421_ (.A(_183_),
    .B(_184_),
    .X(_185_));
 sky130_fd_sc_hd__a22o_1 _422_ (.A1(_097_),
    .A2(net14),
    .B1(_265_),
    .B2(_101_),
    .X(_186_));
 sky130_fd_sc_hd__or3_1 _423_ (.A(_061_),
    .B(_042_),
    .C(_154_),
    .X(_187_));
 sky130_fd_sc_hd__o2111a_1 _424_ (.A1(_266_),
    .A2(_097_),
    .B1(net14),
    .C1(_265_),
    .D1(_301_),
    .X(_188_));
 sky130_fd_sc_hd__and3_1 _425_ (.A(_186_),
    .B(_187_),
    .C(_188_),
    .X(_189_));
 sky130_fd_sc_hd__a21oi_1 _426_ (.A1(_186_),
    .A2(_187_),
    .B1(_188_),
    .Y(_190_));
 sky130_fd_sc_hd__or2_1 _427_ (.A(_189_),
    .B(_190_),
    .X(_191_));
 sky130_fd_sc_hd__xnor2_1 _428_ (.A(_185_),
    .B(_191_),
    .Y(_192_));
 sky130_fd_sc_hd__or2_1 _429_ (.A(_158_),
    .B(_192_),
    .X(_193_));
 sky130_fd_sc_hd__nand2_1 _430_ (.A(_158_),
    .B(_192_),
    .Y(_194_));
 sky130_fd_sc_hd__and2_1 _431_ (.A(_193_),
    .B(_194_),
    .X(_195_));
 sky130_fd_sc_hd__and3_1 _432_ (.A(_121_),
    .B(_162_),
    .C(_164_),
    .X(_196_));
 sky130_fd_sc_hd__xnor2_1 _433_ (.A(_195_),
    .B(_196_),
    .Y(_197_));
 sky130_fd_sc_hd__o21ai_1 _434_ (.A1(_182_),
    .A2(_168_),
    .B1(_197_),
    .Y(_198_));
 sky130_fd_sc_hd__or3_1 _435_ (.A(_182_),
    .B(_168_),
    .C(_197_),
    .X(_199_));
 sky130_fd_sc_hd__and2_1 _436_ (.A(_198_),
    .B(_199_),
    .X(_200_));
 sky130_fd_sc_hd__nand2_1 _437_ (.A(_171_),
    .B(_177_),
    .Y(_201_));
 sky130_fd_sc_hd__a21boi_1 _438_ (.A1(_141_),
    .A2(_172_),
    .B1_N(_139_),
    .Y(_202_));
 sky130_fd_sc_hd__and3_1 _439_ (.A(_175_),
    .B(_201_),
    .C(_202_),
    .X(_203_));
 sky130_fd_sc_hd__xnor2_1 _440_ (.A(_200_),
    .B(_203_),
    .Y(_204_));
 sky130_fd_sc_hd__xor2_1 _441_ (.A(_181_),
    .B(_204_),
    .X(net19));
 sky130_fd_sc_hd__and2b_1 _442_ (.A_N(_203_),
    .B(_200_),
    .X(_205_));
 sky130_fd_sc_hd__a21o_1 _443_ (.A1(_181_),
    .A2(_204_),
    .B1(_205_),
    .X(_206_));
 sky130_fd_sc_hd__or2b_1 _444_ (.A(_196_),
    .B_N(_195_),
    .X(_207_));
 sky130_fd_sc_hd__or2_1 _445_ (.A(_185_),
    .B(_191_),
    .X(_208_));
 sky130_fd_sc_hd__nand2_1 _446_ (.A(_097_),
    .B(_038_),
    .Y(_209_));
 sky130_fd_sc_hd__and3_1 _447_ (.A(_301_),
    .B(_037_),
    .C(_157_),
    .X(_210_));
 sky130_fd_sc_hd__xor2_1 _448_ (.A(_209_),
    .B(_210_),
    .X(_211_));
 sky130_fd_sc_hd__and3_1 _449_ (.A(_101_),
    .B(net14),
    .C(_154_),
    .X(_212_));
 sky130_fd_sc_hd__xnor2_1 _450_ (.A(_189_),
    .B(_212_),
    .Y(_213_));
 sky130_fd_sc_hd__nor2_1 _451_ (.A(_211_),
    .B(_213_),
    .Y(_214_));
 sky130_fd_sc_hd__and2_1 _452_ (.A(_211_),
    .B(_213_),
    .X(_215_));
 sky130_fd_sc_hd__or2_1 _453_ (.A(_214_),
    .B(_215_),
    .X(_216_));
 sky130_fd_sc_hd__a21oi_1 _454_ (.A1(_208_),
    .A2(_193_),
    .B1(_216_),
    .Y(_217_));
 sky130_fd_sc_hd__and3_1 _455_ (.A(_208_),
    .B(_193_),
    .C(_216_),
    .X(_218_));
 sky130_fd_sc_hd__or2_1 _456_ (.A(_217_),
    .B(_218_),
    .X(_219_));
 sky130_fd_sc_hd__a21oi_1 _457_ (.A1(_207_),
    .A2(_198_),
    .B1(_219_),
    .Y(_220_));
 sky130_fd_sc_hd__and3_1 _458_ (.A(_207_),
    .B(_198_),
    .C(_219_),
    .X(_221_));
 sky130_fd_sc_hd__nor2_1 _459_ (.A(_220_),
    .B(_221_),
    .Y(_222_));
 sky130_fd_sc_hd__xor2_1 _460_ (.A(_206_),
    .B(_222_),
    .X(net20));
 sky130_fd_sc_hd__a21bo_1 _461_ (.A1(_189_),
    .A2(_212_),
    .B1_N(_187_),
    .X(_223_));
 sky130_fd_sc_hd__a22o_1 _462_ (.A1(_097_),
    .A2(_037_),
    .B1(_038_),
    .B2(_101_),
    .X(_224_));
 sky130_fd_sc_hd__nand4_1 _463_ (.A(_097_),
    .B(_101_),
    .C(_037_),
    .D(_038_),
    .Y(_225_));
 sky130_fd_sc_hd__a31o_1 _464_ (.A1(_097_),
    .A2(_038_),
    .A3(_210_),
    .B1(_184_),
    .X(_226_));
 sky130_fd_sc_hd__and3_1 _465_ (.A(_224_),
    .B(_225_),
    .C(_226_),
    .X(_228_));
 sky130_fd_sc_hd__a21oi_1 _466_ (.A1(_224_),
    .A2(_225_),
    .B1(_226_),
    .Y(_229_));
 sky130_fd_sc_hd__or2_1 _467_ (.A(_228_),
    .B(_229_),
    .X(_230_));
 sky130_fd_sc_hd__xnor2_1 _468_ (.A(_223_),
    .B(_230_),
    .Y(_231_));
 sky130_fd_sc_hd__o21ai_1 _469_ (.A1(_214_),
    .A2(_217_),
    .B1(_231_),
    .Y(_232_));
 sky130_fd_sc_hd__or3_1 _470_ (.A(_214_),
    .B(_217_),
    .C(_231_),
    .X(_233_));
 sky130_fd_sc_hd__and2_1 _471_ (.A(_232_),
    .B(_233_),
    .X(_234_));
 sky130_fd_sc_hd__a21oi_1 _472_ (.A1(_206_),
    .A2(_222_),
    .B1(_220_),
    .Y(_235_));
 sky130_fd_sc_hd__xnor2_1 _473_ (.A(_234_),
    .B(_235_),
    .Y(net21));
 sky130_fd_sc_hd__and3_1 _474_ (.A(_206_),
    .B(_222_),
    .C(_234_),
    .X(_236_));
 sky130_fd_sc_hd__or2b_1 _475_ (.A(_230_),
    .B_N(_223_),
    .X(_237_));
 sky130_fd_sc_hd__and3_1 _476_ (.A(_101_),
    .B(_037_),
    .C(_209_),
    .X(_238_));
 sky130_fd_sc_hd__nor2_1 _477_ (.A(_228_),
    .B(_238_),
    .Y(_239_));
 sky130_fd_sc_hd__a31o_1 _478_ (.A1(_101_),
    .A2(_037_),
    .A3(_228_),
    .B1(_239_),
    .X(_240_));
 sky130_fd_sc_hd__a21oi_1 _479_ (.A1(_237_),
    .A2(_232_),
    .B1(_240_),
    .Y(_241_));
 sky130_fd_sc_hd__and3_1 _480_ (.A(_237_),
    .B(_232_),
    .C(_240_),
    .X(_242_));
 sky130_fd_sc_hd__nor2_1 _481_ (.A(_241_),
    .B(_242_),
    .Y(_243_));
 sky130_fd_sc_hd__and3_1 _482_ (.A(_220_),
    .B(_234_),
    .C(_243_),
    .X(_244_));
 sky130_fd_sc_hd__a21oi_1 _483_ (.A1(_220_),
    .A2(_234_),
    .B1(_243_),
    .Y(_245_));
 sky130_fd_sc_hd__nor2_1 _484_ (.A(_244_),
    .B(_245_),
    .Y(_246_));
 sky130_fd_sc_hd__xor2_1 _485_ (.A(_236_),
    .B(_246_),
    .X(net22));
 sky130_fd_sc_hd__a21bo_1 _486_ (.A1(_228_),
    .A2(_238_),
    .B1_N(_225_),
    .X(_248_));
 sky130_fd_sc_hd__or2_1 _487_ (.A(_241_),
    .B(_244_),
    .X(_249_));
 sky130_fd_sc_hd__a211o_1 _488_ (.A1(_236_),
    .A2(_246_),
    .B1(_248_),
    .C1(_249_),
    .X(net23));
 sky130_fd_sc_hd__xnor2_1 _489_ (.A(_292_),
    .B(_007_),
    .Y(net28));
 sky130_fd_sc_hd__xor2_1 _490_ (.A(_009_),
    .B(_034_),
    .X(net29));
 sky130_fd_sc_hd__xor2_1 _491_ (.A(_036_),
    .B(_073_),
    .X(net30));
 sky130_fd_sc_hd__xor2_1 _492_ (.A(_075_),
    .B(_111_),
    .X(net31));
 sky130_fd_sc_hd__xor2_1 _493_ (.A(_113_),
    .B(_150_),
    .X(net32));
 sky130_fd_sc_hd__a21oi_1 _494_ (.A1(_253_),
    .A2(_265_),
    .B1(_291_),
    .Y(_250_));
 sky130_fd_sc_hd__nor2_1 _495_ (.A(_292_),
    .B(_250_),
    .Y(net27));
 sky130_fd_sc_hd__or2b_1 _496_ (.A(_279_),
    .B_N(_278_),
    .X(_252_));
 sky130_fd_sc_hd__xnor2_1 _497_ (.A(_264_),
    .B(_252_),
    .Y(net26));
 sky130_fd_sc_hd__nand2_1 _498_ (.A(net1),
    .B(net9),
    .Y(_227_));
 sky130_fd_sc_hd__inv_2 _499_ (.A(_227_),
    .Y(net17));
 sky130_fd_sc_hd__buf_2 _500_ (.A(net10),
    .X(_247_));
 sky130_fd_sc_hd__nand2_1 _501_ (.A(_247_),
    .B(net2),
    .Y(_251_));
 sky130_fd_sc_hd__buf_2 _502_ (.A(net1),
    .X(_253_));
 sky130_fd_sc_hd__buf_2 _503_ (.A(net2),
    .X(_254_));
 sky130_fd_sc_hd__buf_2 _504_ (.A(net9),
    .X(_255_));
 sky130_fd_sc_hd__a22o_1 _505_ (.A1(_253_),
    .A2(_247_),
    .B1(_254_),
    .B2(_255_),
    .X(_256_));
 sky130_fd_sc_hd__o21a_1 _506_ (.A1(_227_),
    .A2(_251_),
    .B1(_256_),
    .X(net24));
 sky130_fd_sc_hd__buf_2 _507_ (.A(net3),
    .X(_257_));
 sky130_fd_sc_hd__nand2_1 _508_ (.A(_255_),
    .B(_257_),
    .Y(_258_));
 sky130_fd_sc_hd__or3b_1 _509_ (.A(_251_),
    .B(_258_),
    .C_N(_227_),
    .X(_259_));
 sky130_fd_sc_hd__a32o_1 _510_ (.A1(_247_),
    .A2(_254_),
    .A3(_227_),
    .B1(_257_),
    .B2(_255_),
    .X(_260_));
 sky130_fd_sc_hd__buf_2 _511_ (.A(net11),
    .X(_261_));
 sky130_fd_sc_hd__and2_1 _512_ (.A(_253_),
    .B(_261_),
    .X(_262_));
 sky130_fd_sc_hd__a21oi_1 _513_ (.A1(_259_),
    .A2(_260_),
    .B1(_262_),
    .Y(_263_));
 sky130_fd_sc_hd__and3_1 _514_ (.A(_259_),
    .B(_260_),
    .C(_262_),
    .X(_264_));
 sky130_fd_sc_hd__nor2_1 _515_ (.A(_263_),
    .B(_264_),
    .Y(net25));
 sky130_fd_sc_hd__buf_2 _516_ (.A(net13),
    .X(_265_));
 sky130_fd_sc_hd__buf_2 _517_ (.A(net5),
    .X(_266_));
 sky130_fd_sc_hd__nand2_1 _518_ (.A(net1),
    .B(_261_),
    .Y(_267_));
 sky130_fd_sc_hd__nand2_1 _519_ (.A(net2),
    .B(net12),
    .Y(_268_));
 sky130_fd_sc_hd__or2_1 _520_ (.A(_267_),
    .B(_268_),
    .X(_269_));
 sky130_fd_sc_hd__clkbuf_2 _521_ (.A(net12),
    .X(_270_));
 sky130_fd_sc_hd__a22o_1 _522_ (.A1(_254_),
    .A2(_261_),
    .B1(_270_),
    .B2(_253_),
    .X(_271_));
 sky130_fd_sc_hd__buf_2 _523_ (.A(net4),
    .X(_272_));
 sky130_fd_sc_hd__nand4_1 _524_ (.A(_255_),
    .B(net10),
    .C(net3),
    .D(_272_),
    .Y(_273_));
 sky130_fd_sc_hd__a22o_1 _525_ (.A1(net10),
    .A2(net3),
    .B1(net4),
    .B2(net9),
    .X(_274_));
 sky130_fd_sc_hd__o2111a_1 _526_ (.A1(net1),
    .A2(net3),
    .B1(net2),
    .C1(net10),
    .D1(net9),
    .X(_275_));
 sky130_fd_sc_hd__a21o_1 _527_ (.A1(_273_),
    .A2(_274_),
    .B1(_275_),
    .X(_276_));
 sky130_fd_sc_hd__nand3_1 _528_ (.A(_273_),
    .B(_274_),
    .C(_275_),
    .Y(_277_));
 sky130_fd_sc_hd__a22o_1 _529_ (.A1(_269_),
    .A2(_271_),
    .B1(_276_),
    .B2(_277_),
    .X(_278_));
 sky130_fd_sc_hd__and4_1 _530_ (.A(_277_),
    .B(_269_),
    .C(_271_),
    .D(_276_),
    .X(_279_));
 sky130_fd_sc_hd__a21o_1 _531_ (.A1(_264_),
    .A2(_278_),
    .B1(_279_),
    .X(_280_));
 sky130_fd_sc_hd__nand2_1 _532_ (.A(net3),
    .B(net11),
    .Y(_281_));
 sky130_fd_sc_hd__nor2_1 _533_ (.A(_262_),
    .B(_268_),
    .Y(_282_));
 sky130_fd_sc_hd__xor2_1 _534_ (.A(_281_),
    .B(_282_),
    .X(_283_));
 sky130_fd_sc_hd__and3_1 _535_ (.A(_273_),
    .B(_274_),
    .C(_275_),
    .X(_284_));
 sky130_fd_sc_hd__and3_1 _536_ (.A(_247_),
    .B(_272_),
    .C(_258_),
    .X(_285_));
 sky130_fd_sc_hd__xnor2_1 _537_ (.A(_284_),
    .B(_285_),
    .Y(_286_));
 sky130_fd_sc_hd__xnor2_1 _538_ (.A(_283_),
    .B(_286_),
    .Y(_287_));
 sky130_fd_sc_hd__xnor2_1 _539_ (.A(_280_),
    .B(_287_),
    .Y(_288_));
 sky130_fd_sc_hd__and3_1 _540_ (.A(_255_),
    .B(_266_),
    .C(_288_),
    .X(_289_));
 sky130_fd_sc_hd__a21oi_1 _541_ (.A1(_255_),
    .A2(_266_),
    .B1(_288_),
    .Y(_290_));
 sky130_fd_sc_hd__nor2_1 _542_ (.A(_289_),
    .B(_290_),
    .Y(_291_));
 sky130_fd_sc_hd__and3_1 _543_ (.A(_253_),
    .B(_265_),
    .C(_291_),
    .X(_292_));
 sky130_fd_sc_hd__inv_2 _544_ (.A(_292_),
    .Y(_293_));
 sky130_fd_sc_hd__nand2_1 _545_ (.A(_253_),
    .B(_265_),
    .Y(_294_));
 sky130_fd_sc_hd__nand2_1 _546_ (.A(_254_),
    .B(net14),
    .Y(_295_));
 sky130_fd_sc_hd__a22o_1 _547_ (.A1(_253_),
    .A2(net14),
    .B1(_265_),
    .B2(_254_),
    .X(_296_));
 sky130_fd_sc_hd__o21ai_2 _548_ (.A1(_294_),
    .A2(_295_),
    .B1(_296_),
    .Y(_297_));
 sky130_fd_sc_hd__inv_2 _549_ (.A(_289_),
    .Y(_298_));
 sky130_fd_sc_hd__nand2_1 _550_ (.A(_255_),
    .B(net5),
    .Y(_299_));
 sky130_fd_sc_hd__nand2_1 _551_ (.A(_247_),
    .B(net6),
    .Y(_300_));
 sky130_fd_sc_hd__buf_2 _552_ (.A(net6),
    .X(_301_));
 sky130_fd_sc_hd__a22o_1 _553_ (.A1(_255_),
    .A2(_301_),
    .B1(_266_),
    .B2(_247_),
    .X(_302_));
 sky130_fd_sc_hd__o21ai_1 _554_ (.A1(_299_),
    .A2(_300_),
    .B1(_302_),
    .Y(_303_));
 sky130_fd_sc_hd__nand2_1 _555_ (.A(_283_),
    .B(_286_),
    .Y(_304_));
 sky130_fd_sc_hd__nor2_1 _556_ (.A(_283_),
    .B(_286_),
    .Y(_305_));
 sky130_fd_sc_hd__a21o_1 _557_ (.A1(_280_),
    .A2(_304_),
    .B1(_305_),
    .X(_306_));
 sky130_fd_sc_hd__a21boi_1 _558_ (.A1(_284_),
    .A2(_285_),
    .B1_N(_273_),
    .Y(_307_));
 sky130_fd_sc_hd__inv_2 _559_ (.A(net4),
    .Y(_308_));
 sky130_fd_sc_hd__inv_2 _560_ (.A(net12),
    .Y(_309_));
 sky130_fd_sc_hd__or3_1 _561_ (.A(_308_),
    .B(_309_),
    .C(_281_),
    .X(_310_));
 sky130_fd_sc_hd__a22o_1 _562_ (.A1(_261_),
    .A2(_272_),
    .B1(net12),
    .B2(_257_),
    .X(_311_));
 sky130_fd_sc_hd__a21oi_1 _563_ (.A1(_267_),
    .A2(_281_),
    .B1(_268_),
    .Y(_312_));
 sky130_fd_sc_hd__and3_1 _564_ (.A(_310_),
    .B(_311_),
    .C(_312_),
    .X(_313_));
 sky130_fd_sc_hd__a21oi_1 _565_ (.A1(_310_),
    .A2(_311_),
    .B1(_312_),
    .Y(_000_));
 sky130_fd_sc_hd__or3_1 _566_ (.A(_307_),
    .B(_313_),
    .C(_000_),
    .X(_001_));
 sky130_fd_sc_hd__o21ai_1 _567_ (.A1(_313_),
    .A2(_000_),
    .B1(_307_),
    .Y(_002_));
 sky130_fd_sc_hd__and2_1 _568_ (.A(_001_),
    .B(_002_),
    .X(_003_));
 sky130_fd_sc_hd__xor2_1 _569_ (.A(_306_),
    .B(_003_),
    .X(_004_));
 sky130_fd_sc_hd__xor2_1 _570_ (.A(_303_),
    .B(_004_),
    .X(_005_));
 sky130_fd_sc_hd__xnor2_1 _571_ (.A(_298_),
    .B(_005_),
    .Y(_006_));
 sky130_fd_sc_hd__xnor2_1 _572_ (.A(_297_),
    .B(_006_),
    .Y(_007_));
 sky130_fd_sc_hd__nor2_1 _573_ (.A(_297_),
    .B(_006_),
    .Y(_008_));
 sky130_fd_sc_hd__o21bai_1 _574_ (.A1(_293_),
    .A2(_007_),
    .B1_N(_008_),
    .Y(_009_));
 sky130_fd_sc_hd__and2_1 _575_ (.A(_253_),
    .B(net15),
    .X(_010_));
 sky130_fd_sc_hd__nand2_1 _576_ (.A(_257_),
    .B(net13),
    .Y(_011_));
 sky130_fd_sc_hd__and3_1 _577_ (.A(_254_),
    .B(net14),
    .C(_294_),
    .X(_012_));
 sky130_fd_sc_hd__xnor2_1 _578_ (.A(_011_),
    .B(_012_),
    .Y(_013_));
 sky130_fd_sc_hd__nand2_1 _579_ (.A(_010_),
    .B(_013_),
    .Y(_014_));
 sky130_fd_sc_hd__or2_1 _580_ (.A(_010_),
    .B(_013_),
    .X(_015_));
 sky130_fd_sc_hd__and2_1 _581_ (.A(_014_),
    .B(_015_),
    .X(_016_));
 sky130_fd_sc_hd__or2b_1 _582_ (.A(_303_),
    .B_N(_004_),
    .X(_017_));
 sky130_fd_sc_hd__o21ai_1 _583_ (.A1(_298_),
    .A2(_005_),
    .B1(_017_),
    .Y(_018_));
 sky130_fd_sc_hd__nand2_1 _584_ (.A(_255_),
    .B(net7),
    .Y(_019_));
 sky130_fd_sc_hd__and3_1 _585_ (.A(_247_),
    .B(net6),
    .C(_299_),
    .X(_020_));
 sky130_fd_sc_hd__xnor2_1 _586_ (.A(_019_),
    .B(_020_),
    .Y(_021_));
 sky130_fd_sc_hd__nand2_1 _587_ (.A(_261_),
    .B(net5),
    .Y(_022_));
 sky130_fd_sc_hd__inv_2 _588_ (.A(_022_),
    .Y(_023_));
 sky130_fd_sc_hd__and2_1 _589_ (.A(_021_),
    .B(_023_),
    .X(_024_));
 sky130_fd_sc_hd__nor2_1 _590_ (.A(_021_),
    .B(_023_),
    .Y(_025_));
 sky130_fd_sc_hd__or2_1 _591_ (.A(_024_),
    .B(_025_),
    .X(_026_));
 sky130_fd_sc_hd__a21bo_1 _592_ (.A1(_306_),
    .A2(_003_),
    .B1_N(_001_),
    .X(_027_));
 sky130_fd_sc_hd__and3_1 _593_ (.A(_272_),
    .B(_270_),
    .C(_313_),
    .X(_028_));
 sky130_fd_sc_hd__a31o_1 _594_ (.A1(_272_),
    .A2(_270_),
    .A3(_281_),
    .B1(_313_),
    .X(_029_));
 sky130_fd_sc_hd__or2b_1 _595_ (.A(_028_),
    .B_N(_029_),
    .X(_030_));
 sky130_fd_sc_hd__xor2_1 _596_ (.A(_027_),
    .B(_030_),
    .X(_031_));
 sky130_fd_sc_hd__xor2_1 _597_ (.A(_026_),
    .B(_031_),
    .X(_032_));
 sky130_fd_sc_hd__xor2_1 _598_ (.A(_018_),
    .B(_032_),
    .X(_033_));
 sky130_fd_sc_hd__xor2_1 _599_ (.A(_016_),
    .B(_033_),
    .X(_034_));
 sky130_fd_sc_hd__and2_1 _600_ (.A(_016_),
    .B(_033_),
    .X(_035_));
 sky130_fd_sc_hd__a21o_1 _601_ (.A1(_009_),
    .A2(_034_),
    .B1(_035_),
    .X(_036_));
 sky130_fd_sc_hd__buf_2 _602_ (.A(net16),
    .X(_037_));
 sky130_fd_sc_hd__buf_2 _603_ (.A(net15),
    .X(_038_));
 sky130_fd_sc_hd__a22oi_1 _604_ (.A1(_253_),
    .A2(net16),
    .B1(_038_),
    .B2(_254_),
    .Y(_039_));
 sky130_fd_sc_hd__a31o_1 _605_ (.A1(_254_),
    .A2(_037_),
    .A3(_010_),
    .B1(_039_),
    .X(_040_));
 sky130_fd_sc_hd__a21oi_1 _606_ (.A1(_011_),
    .A2(_294_),
    .B1(_295_),
    .Y(_041_));
 sky130_fd_sc_hd__inv_2 _607_ (.A(net14),
    .Y(_042_));
 sky130_fd_sc_hd__a22o_1 _608_ (.A1(_257_),
    .A2(net14),
    .B1(net13),
    .B2(_272_),
    .X(_043_));
 sky130_fd_sc_hd__o31a_1 _609_ (.A1(_308_),
    .A2(_042_),
    .A3(_011_),
    .B1(_043_),
    .X(_044_));
 sky130_fd_sc_hd__and2_1 _610_ (.A(_041_),
    .B(_044_),
    .X(_045_));
 sky130_fd_sc_hd__nor2_1 _611_ (.A(_041_),
    .B(_044_),
    .Y(_046_));
 sky130_fd_sc_hd__nor2_1 _612_ (.A(_045_),
    .B(_046_),
    .Y(_047_));
 sky130_fd_sc_hd__xor2_1 _613_ (.A(_040_),
    .B(_047_),
    .X(_048_));
 sky130_fd_sc_hd__nor2_1 _614_ (.A(_014_),
    .B(_048_),
    .Y(_049_));
 sky130_fd_sc_hd__and2_1 _615_ (.A(_014_),
    .B(_048_),
    .X(_050_));
 sky130_fd_sc_hd__nor2_1 _616_ (.A(_049_),
    .B(_050_),
    .Y(_051_));
 sky130_fd_sc_hd__nor2_1 _617_ (.A(_026_),
    .B(_031_),
    .Y(_052_));
 sky130_fd_sc_hd__a21o_1 _618_ (.A1(_018_),
    .A2(_032_),
    .B1(_052_),
    .X(_053_));
 sky130_fd_sc_hd__and4_1 _619_ (.A(_257_),
    .B(_261_),
    .C(_272_),
    .D(_270_),
    .X(_054_));
 sky130_fd_sc_hd__and2b_1 _620_ (.A_N(_030_),
    .B(_027_),
    .X(_055_));
 sky130_fd_sc_hd__a22oi_1 _621_ (.A1(_261_),
    .A2(_301_),
    .B1(_266_),
    .B2(_270_),
    .Y(_056_));
 sky130_fd_sc_hd__and3_1 _622_ (.A(_270_),
    .B(net6),
    .C(_023_),
    .X(_057_));
 sky130_fd_sc_hd__or2_1 _623_ (.A(_056_),
    .B(_057_),
    .X(_058_));
 sky130_fd_sc_hd__a22o_1 _624_ (.A1(_247_),
    .A2(net7),
    .B1(net8),
    .B2(_255_),
    .X(_059_));
 sky130_fd_sc_hd__inv_2 _625_ (.A(_247_),
    .Y(_060_));
 sky130_fd_sc_hd__inv_2 _626_ (.A(net8),
    .Y(_061_));
 sky130_fd_sc_hd__or3_1 _627_ (.A(_060_),
    .B(_061_),
    .C(_019_),
    .X(_062_));
 sky130_fd_sc_hd__a21oi_1 _628_ (.A1(_019_),
    .A2(_299_),
    .B1(_300_),
    .Y(_063_));
 sky130_fd_sc_hd__and3_1 _629_ (.A(_059_),
    .B(_062_),
    .C(_063_),
    .X(_064_));
 sky130_fd_sc_hd__a21oi_1 _630_ (.A1(_059_),
    .A2(_062_),
    .B1(_063_),
    .Y(_065_));
 sky130_fd_sc_hd__or2_1 _631_ (.A(_064_),
    .B(_065_),
    .X(_066_));
 sky130_fd_sc_hd__xnor2_1 _632_ (.A(_058_),
    .B(_066_),
    .Y(_067_));
 sky130_fd_sc_hd__xnor2_1 _633_ (.A(_024_),
    .B(_067_),
    .Y(_068_));
 sky130_fd_sc_hd__o31a_1 _634_ (.A1(_054_),
    .A2(_028_),
    .A3(_055_),
    .B1(_068_),
    .X(_069_));
 sky130_fd_sc_hd__or4_1 _635_ (.A(_068_),
    .B(_054_),
    .C(_028_),
    .D(_055_),
    .X(_070_));
 sky130_fd_sc_hd__or2b_1 _636_ (.A(_069_),
    .B_N(_070_),
    .X(_071_));
 sky130_fd_sc_hd__xnor2_1 _637_ (.A(_053_),
    .B(_071_),
    .Y(_072_));
 sky130_fd_sc_hd__xor2_1 _638_ (.A(_051_),
    .B(_072_),
    .X(_073_));
 sky130_fd_sc_hd__and2_1 _639_ (.A(_051_),
    .B(_072_),
    .X(_074_));
 sky130_fd_sc_hd__a21o_1 _640_ (.A1(_036_),
    .A2(_073_),
    .B1(_074_),
    .X(_075_));
 sky130_fd_sc_hd__and2b_1 _641_ (.A_N(_040_),
    .B(_047_),
    .X(_076_));
 sky130_fd_sc_hd__nand2_1 _642_ (.A(_257_),
    .B(net15),
    .Y(_077_));
 sky130_fd_sc_hd__and3b_1 _643_ (.A_N(_010_),
    .B(net16),
    .C(_254_),
    .X(_078_));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_130 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(a[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(a[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(a[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(a[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(a[4]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(a[5]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(a[6]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(a[7]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(b[0]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(b[1]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(b[2]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(b[3]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(b[4]),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input14 (.A(b[5]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(b[6]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(b[7]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(prod[0]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(prod[10]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(prod[11]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(prod[12]));
 sky130_fd_sc_hd__clkbuf_4 output21 (.A(net21),
    .X(prod[13]));
 sky130_fd_sc_hd__clkbuf_4 output22 (.A(net22),
    .X(prod[14]));
 sky130_fd_sc_hd__clkbuf_4 output23 (.A(net23),
    .X(prod[15]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(prod[1]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(prod[2]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(prod[3]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(prod[4]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(prod[5]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(prod[6]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(prod[7]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(prod[8]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(prod[9]));
endmodule
