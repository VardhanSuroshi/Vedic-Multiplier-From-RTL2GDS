VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pes_vedic_mul
  CLASS BLOCK ;
  FOREIGN pes_vedic_mul ;
  ORIGIN 0.000 0.000 ;
  SIZE 87.495 BY 98.215 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 17.565 10.640 19.165 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.655 10.640 38.255 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 55.745 10.640 57.345 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.835 10.640 76.435 87.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 22.900 82.120 24.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 41.940 82.120 43.540 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 60.980 82.120 62.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 80.020 82.120 81.620 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.265 10.640 15.865 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 33.355 10.640 34.955 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 52.445 10.640 54.045 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.535 10.640 73.135 87.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 19.600 82.120 21.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 38.640 82.120 40.240 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 57.680 82.120 59.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 76.720 82.120 78.320 ;
    END
  END VPWR
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END a[0]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END a[7]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END b[0]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END b[1]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END b[2]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END b[3]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END b[4]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END b[5]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END b[7]
  PIN prod[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END prod[0]
  PIN prod[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 83.495 54.440 87.495 55.040 ;
    END
  END prod[10]
  PIN prod[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 83.495 64.640 87.495 65.240 ;
    END
  END prod[11]
  PIN prod[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 83.495 74.840 87.495 75.440 ;
    END
  END prod[12]
  PIN prod[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 74.150 94.215 74.430 98.215 ;
    END
  END prod[13]
  PIN prod[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 67.710 94.215 67.990 98.215 ;
    END
  END prod[14]
  PIN prod[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 94.215 61.550 98.215 ;
    END
  END prod[15]
  PIN prod[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END prod[1]
  PIN prod[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END prod[2]
  PIN prod[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END prod[3]
  PIN prod[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END prod[4]
  PIN prod[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END prod[5]
  PIN prod[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 83.495 17.040 87.495 17.640 ;
    END
  END prod[6]
  PIN prod[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 83.495 27.240 87.495 27.840 ;
    END
  END prod[7]
  PIN prod[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 83.495 37.440 87.495 38.040 ;
    END
  END prod[8]
  PIN prod[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 83.495 47.640 87.495 48.240 ;
    END
  END prod[9]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 81.880 87.125 ;
      LAYER met1 ;
        RECT 4.670 10.640 81.880 87.280 ;
      LAYER met2 ;
        RECT 4.690 93.935 60.990 94.930 ;
        RECT 61.830 93.935 67.430 94.930 ;
        RECT 68.270 93.935 73.870 94.930 ;
        RECT 74.710 93.935 80.410 94.930 ;
        RECT 4.690 4.280 80.410 93.935 ;
        RECT 4.690 4.000 22.350 4.280 ;
        RECT 23.190 4.000 35.230 4.280 ;
        RECT 36.070 4.000 38.450 4.280 ;
        RECT 39.290 4.000 41.670 4.280 ;
        RECT 42.510 4.000 44.890 4.280 ;
        RECT 45.730 4.000 60.990 4.280 ;
        RECT 61.830 4.000 80.410 4.280 ;
      LAYER met3 ;
        RECT 4.000 75.840 83.495 87.205 ;
        RECT 4.000 74.440 83.095 75.840 ;
        RECT 4.000 72.440 83.495 74.440 ;
        RECT 4.400 71.040 83.495 72.440 ;
        RECT 4.000 65.640 83.495 71.040 ;
        RECT 4.400 64.240 83.095 65.640 ;
        RECT 4.000 62.240 83.495 64.240 ;
        RECT 4.400 60.840 83.495 62.240 ;
        RECT 4.000 55.440 83.495 60.840 ;
        RECT 4.400 54.040 83.095 55.440 ;
        RECT 4.000 52.040 83.495 54.040 ;
        RECT 4.400 50.640 83.495 52.040 ;
        RECT 4.000 48.640 83.495 50.640 ;
        RECT 4.400 47.240 83.095 48.640 ;
        RECT 4.000 45.240 83.495 47.240 ;
        RECT 4.400 43.840 83.495 45.240 ;
        RECT 4.000 41.840 83.495 43.840 ;
        RECT 4.400 40.440 83.495 41.840 ;
        RECT 4.000 38.440 83.495 40.440 ;
        RECT 4.400 37.040 83.095 38.440 ;
        RECT 4.000 35.040 83.495 37.040 ;
        RECT 4.400 33.640 83.495 35.040 ;
        RECT 4.000 31.640 83.495 33.640 ;
        RECT 4.400 30.240 83.495 31.640 ;
        RECT 4.000 28.240 83.495 30.240 ;
        RECT 4.400 26.840 83.095 28.240 ;
        RECT 4.000 24.840 83.495 26.840 ;
        RECT 4.400 23.440 83.495 24.840 ;
        RECT 4.000 21.440 83.495 23.440 ;
        RECT 4.400 20.040 83.495 21.440 ;
        RECT 4.000 18.040 83.495 20.040 ;
        RECT 4.400 16.640 83.095 18.040 ;
        RECT 4.000 14.640 83.495 16.640 ;
        RECT 4.400 13.240 83.495 14.640 ;
        RECT 4.000 10.715 83.495 13.240 ;
  END
END pes_vedic_mul
END LIBRARY

