magic
tech sky130A
magscale 1 2
timestamp 1699032935
<< viali >>
rect 14289 17289 14323 17323
rect 15301 17289 15335 17323
rect 12541 17221 12575 17255
rect 7205 17153 7239 17187
rect 7389 17153 7423 17187
rect 10333 17153 10367 17187
rect 10425 17153 10459 17187
rect 10609 17153 10643 17187
rect 12173 17153 12207 17187
rect 12909 17153 12943 17187
rect 13093 17153 13127 17187
rect 14197 17153 14231 17187
rect 15025 17153 15059 17187
rect 7573 16949 7607 16983
rect 10609 16949 10643 16983
rect 12909 16949 12943 16983
rect 6653 16745 6687 16779
rect 9689 16745 9723 16779
rect 10241 16745 10275 16779
rect 10885 16745 10919 16779
rect 11897 16745 11931 16779
rect 12081 16745 12115 16779
rect 12173 16745 12207 16779
rect 13369 16745 13403 16779
rect 14565 16745 14599 16779
rect 8309 16677 8343 16711
rect 9505 16677 9539 16711
rect 10057 16677 10091 16711
rect 11529 16677 11563 16711
rect 9045 16609 9079 16643
rect 11161 16609 11195 16643
rect 12909 16609 12943 16643
rect 14381 16609 14415 16643
rect 6377 16541 6411 16575
rect 6929 16541 6963 16575
rect 7297 16541 7331 16575
rect 7389 16541 7423 16575
rect 7573 16541 7607 16575
rect 7757 16541 7791 16575
rect 7849 16541 7883 16575
rect 7941 16541 7975 16575
rect 8033 16541 8067 16575
rect 8309 16541 8343 16575
rect 8493 16541 8527 16575
rect 9137 16541 9171 16575
rect 9597 16541 9631 16575
rect 10241 16541 10275 16575
rect 10333 16541 10367 16575
rect 11345 16541 11379 16575
rect 12371 16551 12405 16585
rect 12522 16541 12556 16575
rect 12633 16541 12667 16575
rect 12725 16541 12759 16575
rect 13001 16541 13035 16575
rect 14289 16541 14323 16575
rect 6653 16473 6687 16507
rect 10701 16473 10735 16507
rect 10901 16473 10935 16507
rect 11713 16473 11747 16507
rect 6469 16405 6503 16439
rect 8217 16405 8251 16439
rect 10609 16405 10643 16439
rect 11069 16405 11103 16439
rect 11913 16405 11947 16439
rect 5825 16201 5859 16235
rect 7665 16201 7699 16235
rect 11621 16201 11655 16235
rect 12541 16201 12575 16235
rect 12817 16201 12851 16235
rect 13645 16201 13679 16235
rect 5733 16133 5767 16167
rect 6653 16133 6687 16167
rect 7297 16133 7331 16167
rect 7497 16133 7531 16167
rect 12173 16133 12207 16167
rect 12633 16133 12667 16167
rect 13797 16133 13831 16167
rect 14013 16133 14047 16167
rect 14197 16133 14231 16167
rect 5641 16065 5675 16099
rect 6009 16065 6043 16099
rect 6561 16065 6595 16099
rect 6745 16065 6779 16099
rect 6929 16065 6963 16099
rect 10057 16065 10091 16099
rect 11529 16065 11563 16099
rect 11713 16065 11747 16099
rect 12357 16065 12391 16099
rect 12909 16065 12943 16099
rect 14105 16065 14139 16099
rect 14381 16065 14415 16099
rect 10333 15997 10367 16031
rect 5917 15929 5951 15963
rect 6377 15929 6411 15963
rect 10149 15929 10183 15963
rect 12633 15929 12667 15963
rect 14381 15929 14415 15963
rect 7481 15861 7515 15895
rect 10241 15861 10275 15895
rect 13829 15861 13863 15895
rect 6745 15657 6779 15691
rect 6929 15657 6963 15691
rect 7389 15657 7423 15691
rect 7849 15521 7883 15555
rect 8125 15521 8159 15555
rect 9137 15521 9171 15555
rect 7297 15453 7331 15487
rect 7481 15453 7515 15487
rect 7757 15453 7791 15487
rect 9321 15453 9355 15487
rect 9597 15453 9631 15487
rect 9781 15453 9815 15487
rect 10057 15453 10091 15487
rect 6561 15385 6595 15419
rect 9505 15385 9539 15419
rect 9873 15385 9907 15419
rect 15669 15385 15703 15419
rect 6761 15317 6795 15351
rect 9689 15317 9723 15351
rect 10241 15317 10275 15351
rect 15945 15317 15979 15351
rect 4169 15113 4203 15147
rect 6745 15113 6779 15147
rect 10717 15113 10751 15147
rect 10885 15113 10919 15147
rect 13293 15113 13327 15147
rect 4077 15045 4111 15079
rect 10149 15045 10183 15079
rect 10517 15045 10551 15079
rect 10977 15045 11011 15079
rect 12541 15045 12575 15079
rect 13093 15045 13127 15079
rect 14289 15045 14323 15079
rect 2697 14977 2731 15011
rect 3985 14977 4019 15011
rect 4261 14977 4295 15011
rect 4537 14977 4571 15011
rect 4721 14977 4755 15011
rect 7021 14977 7055 15011
rect 7113 14977 7147 15011
rect 10333 14977 10367 15011
rect 10425 14977 10459 15011
rect 11161 14977 11195 15011
rect 12449 14977 12483 15011
rect 12817 14977 12851 15011
rect 13737 14977 13771 15011
rect 14197 14977 14231 15011
rect 14381 14977 14415 15011
rect 6929 14909 6963 14943
rect 7205 14909 7239 14943
rect 11345 14909 11379 14943
rect 13001 14909 13035 14943
rect 13829 14909 13863 14943
rect 14105 14909 14139 14943
rect 13461 14841 13495 14875
rect 2513 14773 2547 14807
rect 4629 14773 4663 14807
rect 10149 14773 10183 14807
rect 10701 14773 10735 14807
rect 13277 14773 13311 14807
rect 4629 14569 4663 14603
rect 5641 14569 5675 14603
rect 9413 14569 9447 14603
rect 10057 14569 10091 14603
rect 10977 14569 11011 14603
rect 12449 14569 12483 14603
rect 12817 14569 12851 14603
rect 3341 14501 3375 14535
rect 4445 14501 4479 14535
rect 5825 14501 5859 14535
rect 3801 14433 3835 14467
rect 4077 14433 4111 14467
rect 4262 14433 4296 14467
rect 6009 14433 6043 14467
rect 9045 14433 9079 14467
rect 11069 14433 11103 14467
rect 11805 14433 11839 14467
rect 2513 14365 2547 14399
rect 2697 14365 2731 14399
rect 2881 14365 2915 14399
rect 3341 14365 3375 14399
rect 3617 14365 3651 14399
rect 3985 14365 4019 14399
rect 4169 14365 4203 14399
rect 4905 14365 4939 14399
rect 5181 14365 5215 14399
rect 5917 14365 5951 14399
rect 6101 14365 6135 14399
rect 9137 14365 9171 14399
rect 11253 14365 11287 14399
rect 11437 14365 11471 14399
rect 11897 14365 11931 14399
rect 12357 14365 12391 14399
rect 1501 14297 1535 14331
rect 2789 14297 2823 14331
rect 3525 14297 3559 14331
rect 4813 14297 4847 14331
rect 5457 14297 5491 14331
rect 7205 14297 7239 14331
rect 7389 14297 7423 14331
rect 9689 14297 9723 14331
rect 9873 14297 9907 14331
rect 10609 14297 10643 14331
rect 10793 14297 10827 14331
rect 1593 14229 1627 14263
rect 3065 14229 3099 14263
rect 4603 14229 4637 14263
rect 4997 14229 5031 14263
rect 5365 14229 5399 14263
rect 5657 14229 5691 14263
rect 7573 14229 7607 14263
rect 12265 14229 12299 14263
rect 2697 14025 2731 14059
rect 3617 14025 3651 14059
rect 5273 14025 5307 14059
rect 6745 14025 6779 14059
rect 7021 14025 7055 14059
rect 8953 14025 8987 14059
rect 9413 14025 9447 14059
rect 10885 14025 10919 14059
rect 1593 13957 1627 13991
rect 1685 13957 1719 13991
rect 2329 13957 2363 13991
rect 4997 13957 5031 13991
rect 7435 13957 7469 13991
rect 9229 13957 9263 13991
rect 1496 13895 1530 13929
rect 1869 13889 1903 13923
rect 2237 13889 2271 13923
rect 2421 13889 2455 13923
rect 2973 13889 3007 13923
rect 3249 13889 3283 13923
rect 4169 13889 4203 13923
rect 4353 13889 4387 13923
rect 5181 13889 5215 13923
rect 5273 13889 5307 13923
rect 6929 13889 6963 13923
rect 7113 13889 7147 13923
rect 7573 13889 7607 13923
rect 7665 13889 7699 13923
rect 7762 13911 7796 13945
rect 9045 13889 9079 13923
rect 9689 13889 9723 13923
rect 10701 13889 10735 13923
rect 10885 13889 10919 13923
rect 1961 13821 1995 13855
rect 3341 13821 3375 13855
rect 7481 13821 7515 13855
rect 8309 13821 8343 13855
rect 8677 13821 8711 13855
rect 8769 13821 8803 13855
rect 9597 13821 9631 13855
rect 2053 13753 2087 13787
rect 7297 13753 7331 13787
rect 10057 13753 10091 13787
rect 1869 13685 1903 13719
rect 3065 13685 3099 13719
rect 3249 13685 3283 13719
rect 4169 13685 4203 13719
rect 3065 13481 3099 13515
rect 3525 13481 3559 13515
rect 5917 13481 5951 13515
rect 7021 13481 7055 13515
rect 7205 13481 7239 13515
rect 8401 13481 8435 13515
rect 8585 13481 8619 13515
rect 9229 13481 9263 13515
rect 12817 13481 12851 13515
rect 14105 13481 14139 13515
rect 12633 13413 12667 13447
rect 1961 13345 1995 13379
rect 2145 13345 2179 13379
rect 10793 13345 10827 13379
rect 12541 13345 12575 13379
rect 12909 13345 12943 13379
rect 13277 13345 13311 13379
rect 1409 13277 1443 13311
rect 2053 13277 2087 13311
rect 2237 13277 2271 13311
rect 3249 13277 3283 13311
rect 3341 13277 3375 13311
rect 5089 13277 5123 13311
rect 5273 13277 5307 13311
rect 5365 13277 5399 13311
rect 5825 13277 5859 13311
rect 6101 13277 6135 13311
rect 6745 13277 6779 13311
rect 7481 13277 7515 13311
rect 7665 13277 7699 13311
rect 8953 13277 8987 13311
rect 10149 13277 10183 13311
rect 10701 13277 10735 13311
rect 10885 13277 10919 13311
rect 11437 13277 11471 13311
rect 11621 13277 11655 13311
rect 12357 13277 12391 13311
rect 12725 13277 12759 13311
rect 12817 13277 12851 13311
rect 13461 13277 13495 13311
rect 14289 13277 14323 13311
rect 14565 13277 14599 13311
rect 15761 13277 15795 13311
rect 6009 13209 6043 13243
rect 7389 13209 7423 13243
rect 8217 13209 8251 13243
rect 9045 13209 9079 13243
rect 9229 13209 9263 13243
rect 10333 13209 10367 13243
rect 10517 13209 10551 13243
rect 1593 13141 1627 13175
rect 2421 13141 2455 13175
rect 4905 13141 4939 13175
rect 6561 13141 6595 13175
rect 7189 13141 7223 13175
rect 7573 13141 7607 13175
rect 8417 13141 8451 13175
rect 11529 13141 11563 13175
rect 13185 13141 13219 13175
rect 13645 13141 13679 13175
rect 14473 13141 14507 13175
rect 15945 13141 15979 13175
rect 2697 12937 2731 12971
rect 5549 12937 5583 12971
rect 5917 12937 5951 12971
rect 7665 12937 7699 12971
rect 8309 12937 8343 12971
rect 8769 12937 8803 12971
rect 10333 12937 10367 12971
rect 7297 12869 7331 12903
rect 8401 12869 8435 12903
rect 8617 12869 8651 12903
rect 1409 12801 1443 12835
rect 2237 12801 2271 12835
rect 2513 12801 2547 12835
rect 2697 12801 2731 12835
rect 4629 12801 4663 12835
rect 4813 12801 4847 12835
rect 5733 12801 5767 12835
rect 6009 12801 6043 12835
rect 7205 12801 7239 12835
rect 7389 12801 7423 12835
rect 7757 12801 7791 12835
rect 7941 12801 7975 12835
rect 8033 12801 8067 12835
rect 8125 12801 8159 12835
rect 10149 12801 10183 12835
rect 10333 12801 10367 12835
rect 11713 12801 11747 12835
rect 13461 12801 13495 12835
rect 14565 12801 14599 12835
rect 2421 12733 2455 12767
rect 6929 12733 6963 12767
rect 11621 12733 11655 12767
rect 13369 12733 13403 12767
rect 14473 12733 14507 12767
rect 14933 12733 14967 12767
rect 1593 12665 1627 12699
rect 13829 12665 13863 12699
rect 2053 12597 2087 12631
rect 4721 12597 4755 12631
rect 7021 12597 7055 12631
rect 8585 12597 8619 12631
rect 12081 12597 12115 12631
rect 2053 12393 2087 12427
rect 4445 12393 4479 12427
rect 5917 12393 5951 12427
rect 7941 12393 7975 12427
rect 8309 12393 8343 12427
rect 9505 12393 9539 12427
rect 12357 12393 12391 12427
rect 13921 12393 13955 12427
rect 2237 12325 2271 12359
rect 11989 12325 12023 12359
rect 12541 12325 12575 12359
rect 13737 12325 13771 12359
rect 2421 12257 2455 12291
rect 2881 12257 2915 12291
rect 4537 12257 4571 12291
rect 5273 12257 5307 12291
rect 5733 12257 5767 12291
rect 6285 12257 6319 12291
rect 9045 12257 9079 12291
rect 1685 12189 1719 12223
rect 2513 12189 2547 12223
rect 3433 12189 3467 12223
rect 3985 12189 4019 12223
rect 4261 12189 4295 12223
rect 4721 12189 4755 12223
rect 5641 12189 5675 12223
rect 5917 12189 5951 12223
rect 6101 12189 6135 12223
rect 6193 12189 6227 12223
rect 6377 12189 6411 12223
rect 7665 12189 7699 12223
rect 7849 12189 7883 12223
rect 7941 12189 7975 12223
rect 8033 12189 8067 12223
rect 9137 12189 9171 12223
rect 11897 12189 11931 12223
rect 12173 12189 12207 12223
rect 12449 12189 12483 12223
rect 12817 12189 12851 12223
rect 13001 12189 13035 12223
rect 2053 12121 2087 12155
rect 3249 12121 3283 12155
rect 7757 12121 7791 12155
rect 12725 12121 12759 12155
rect 13461 12121 13495 12155
rect 3617 12053 3651 12087
rect 4077 12053 4111 12087
rect 4905 12053 4939 12087
rect 12449 12053 12483 12087
rect 12909 12053 12943 12087
rect 4169 11849 4203 11883
rect 8769 11849 8803 11883
rect 10717 11849 10751 11883
rect 10885 11849 10919 11883
rect 11621 11849 11655 11883
rect 14841 11849 14875 11883
rect 4353 11781 4387 11815
rect 8401 11781 8435 11815
rect 8601 11781 8635 11815
rect 9689 11781 9723 11815
rect 10517 11781 10551 11815
rect 15209 11781 15243 11815
rect 3249 11713 3283 11747
rect 3433 11713 3467 11747
rect 3709 11713 3743 11747
rect 4077 11713 4111 11747
rect 4169 11713 4203 11747
rect 9597 11713 9631 11747
rect 9781 11713 9815 11747
rect 10057 11713 10091 11747
rect 11529 11713 11563 11747
rect 11713 11713 11747 11747
rect 14381 11713 14415 11747
rect 15025 11713 15059 11747
rect 15301 11713 15335 11747
rect 3341 11645 3375 11679
rect 3525 11645 3559 11679
rect 10149 11645 10183 11679
rect 10425 11645 10459 11679
rect 14289 11645 14323 11679
rect 14749 11645 14783 11679
rect 3893 11509 3927 11543
rect 8585 11509 8619 11543
rect 10701 11509 10735 11543
rect 6469 11305 6503 11339
rect 8309 11305 8343 11339
rect 8677 11305 8711 11339
rect 11805 11305 11839 11339
rect 14749 11305 14783 11339
rect 1593 11237 1627 11271
rect 8125 11237 8159 11271
rect 7389 11169 7423 11203
rect 8401 11169 8435 11203
rect 9045 11169 9079 11203
rect 10977 11169 11011 11203
rect 11437 11169 11471 11203
rect 13461 11169 13495 11203
rect 13737 11169 13771 11203
rect 15209 11169 15243 11203
rect 15669 11169 15703 11203
rect 1409 11101 1443 11135
rect 6653 11101 6687 11135
rect 6929 11101 6963 11135
rect 7021 11101 7055 11135
rect 7297 11101 7331 11135
rect 7481 11101 7515 11135
rect 7573 11101 7607 11135
rect 7965 11101 7999 11135
rect 8309 11101 8343 11135
rect 8953 11101 8987 11135
rect 11069 11101 11103 11135
rect 11253 11101 11287 11135
rect 11621 11101 11655 11135
rect 11897 11091 11931 11125
rect 12081 11101 12115 11135
rect 12173 11101 12207 11135
rect 12357 11101 12391 11135
rect 13369 11101 13403 11135
rect 14381 11101 14415 11135
rect 14565 11101 14599 11135
rect 15301 11101 15335 11135
rect 7113 11033 7147 11067
rect 7757 11033 7791 11067
rect 7849 11033 7883 11067
rect 10609 11033 10643 11067
rect 10793 11033 10827 11067
rect 12541 11033 12575 11067
rect 6745 10965 6779 10999
rect 11253 10965 11287 10999
rect 12081 10965 12115 10999
rect 5549 10761 5583 10795
rect 13201 10761 13235 10795
rect 13369 10761 13403 10795
rect 15945 10761 15979 10795
rect 2513 10693 2547 10727
rect 4445 10693 4479 10727
rect 4537 10693 4571 10727
rect 13001 10693 13035 10727
rect 15669 10693 15703 10727
rect 1409 10625 1443 10659
rect 2053 10625 2087 10659
rect 3709 10625 3743 10659
rect 4813 10625 4847 10659
rect 5365 10625 5399 10659
rect 5641 10625 5675 10659
rect 5825 10625 5859 10659
rect 6009 10625 6043 10659
rect 6101 10625 6135 10659
rect 6653 10625 6687 10659
rect 7297 10625 7331 10659
rect 12725 10625 12759 10659
rect 12909 10625 12943 10659
rect 13461 10625 13495 10659
rect 13645 10625 13679 10659
rect 2145 10557 2179 10591
rect 2421 10557 2455 10591
rect 2973 10557 3007 10591
rect 3801 10557 3835 10591
rect 4629 10557 4663 10591
rect 5181 10557 5215 10591
rect 5917 10557 5951 10591
rect 6377 10557 6411 10591
rect 12541 10557 12575 10591
rect 2881 10489 2915 10523
rect 13553 10489 13587 10523
rect 1593 10421 1627 10455
rect 3893 10421 3927 10455
rect 4077 10421 4111 10455
rect 7481 10421 7515 10455
rect 13185 10421 13219 10455
rect 3433 10217 3467 10251
rect 5181 10217 5215 10251
rect 6009 10217 6043 10251
rect 6377 10217 6411 10251
rect 8309 10217 8343 10251
rect 9597 10217 9631 10251
rect 12357 10217 12391 10251
rect 12725 10217 12759 10251
rect 14933 10217 14967 10251
rect 9873 10149 9907 10183
rect 4997 10081 5031 10115
rect 9137 10081 9171 10115
rect 10333 10081 10367 10115
rect 1777 10013 1811 10047
rect 3249 10013 3283 10047
rect 3433 10013 3467 10047
rect 3801 10013 3835 10047
rect 3985 10013 4019 10047
rect 4169 10013 4203 10047
rect 4261 10013 4295 10047
rect 4445 10013 4479 10047
rect 4537 10013 4571 10047
rect 4721 10013 4755 10047
rect 4905 10013 4939 10047
rect 5089 10013 5123 10047
rect 5181 10013 5215 10047
rect 5365 10013 5399 10047
rect 5917 10013 5951 10047
rect 6101 10013 6135 10047
rect 6561 10013 6595 10047
rect 6745 10013 6779 10047
rect 6929 10013 6963 10047
rect 9229 10013 9263 10047
rect 9321 10013 9355 10047
rect 9413 10013 9447 10047
rect 9689 10013 9723 10047
rect 10149 10013 10183 10047
rect 10241 10013 10275 10047
rect 10425 10013 10459 10047
rect 11897 10013 11931 10047
rect 12173 10013 12207 10047
rect 12449 10013 12483 10047
rect 12725 10013 12759 10047
rect 15117 10013 15151 10047
rect 15393 10013 15427 10047
rect 6653 9945 6687 9979
rect 8125 9945 8159 9979
rect 8341 9945 8375 9979
rect 12633 9945 12667 9979
rect 15669 9945 15703 9979
rect 1501 9877 1535 9911
rect 4353 9877 4387 9911
rect 4721 9877 4755 9911
rect 8493 9877 8527 9911
rect 10057 9877 10091 9911
rect 11989 9877 12023 9911
rect 15301 9877 15335 9911
rect 15945 9877 15979 9911
rect 3157 9673 3191 9707
rect 7665 9673 7699 9707
rect 13369 9673 13403 9707
rect 4169 9605 4203 9639
rect 4353 9605 4387 9639
rect 8309 9605 8343 9639
rect 8493 9605 8527 9639
rect 9045 9605 9079 9639
rect 11161 9605 11195 9639
rect 9275 9571 9309 9605
rect 3065 9537 3099 9571
rect 3249 9537 3283 9571
rect 3525 9537 3559 9571
rect 3709 9537 3743 9571
rect 3985 9537 4019 9571
rect 7113 9537 7147 9571
rect 7297 9537 7331 9571
rect 7389 9537 7423 9571
rect 7481 9537 7515 9571
rect 7757 9537 7791 9571
rect 8217 9537 8251 9571
rect 10425 9537 10459 9571
rect 10885 9537 10919 9571
rect 11713 9537 11747 9571
rect 13185 9537 13219 9571
rect 13553 9537 13587 9571
rect 13737 9537 13771 9571
rect 14841 9537 14875 9571
rect 15485 9537 15519 9571
rect 7849 9469 7883 9503
rect 10517 9469 10551 9503
rect 11161 9469 11195 9503
rect 11529 9469 11563 9503
rect 13001 9469 13035 9503
rect 14565 9469 14599 9503
rect 14749 9469 14783 9503
rect 15209 9469 15243 9503
rect 15577 9469 15611 9503
rect 15853 9469 15887 9503
rect 8125 9401 8159 9435
rect 8493 9401 8527 9435
rect 9413 9401 9447 9435
rect 10977 9401 11011 9435
rect 3893 9333 3927 9367
rect 7941 9333 7975 9367
rect 9229 9333 9263 9367
rect 10425 9333 10459 9367
rect 10793 9333 10827 9367
rect 11897 9333 11931 9367
rect 4721 9129 4755 9163
rect 5457 9129 5491 9163
rect 7021 9129 7055 9163
rect 12081 9129 12115 9163
rect 12357 9129 12391 9163
rect 13185 9129 13219 9163
rect 14841 9129 14875 9163
rect 5273 9061 5307 9095
rect 7481 9061 7515 9095
rect 11621 9061 11655 9095
rect 12173 9061 12207 9095
rect 5089 8993 5123 9027
rect 8125 8993 8159 9027
rect 8217 8993 8251 9027
rect 9045 8993 9079 9027
rect 9505 8993 9539 9027
rect 12265 8993 12299 9027
rect 12817 8993 12851 9027
rect 4997 8925 5031 8959
rect 5917 8925 5951 8959
rect 6101 8925 6135 8959
rect 6285 8925 6319 8959
rect 6561 8925 6595 8959
rect 6745 8925 6779 8959
rect 7389 8925 7423 8959
rect 7573 8925 7607 8959
rect 8033 8925 8067 8959
rect 8309 8925 8343 8959
rect 9137 8925 9171 8959
rect 11437 8925 11471 8959
rect 11621 8925 11655 8959
rect 11989 8925 12023 8959
rect 12357 8925 12391 8959
rect 12449 8925 12483 8959
rect 13001 8925 13035 8959
rect 14657 8925 14691 8959
rect 14841 8925 14875 8959
rect 1409 8857 1443 8891
rect 1777 8857 1811 8891
rect 5641 8857 5675 8891
rect 6193 8857 6227 8891
rect 7113 8857 7147 8891
rect 5441 8789 5475 8823
rect 6469 8789 6503 8823
rect 8493 8789 8527 8823
rect 12725 8789 12759 8823
rect 5457 8585 5491 8619
rect 5825 8585 5859 8619
rect 7757 8585 7791 8619
rect 8401 8585 8435 8619
rect 9965 8585 9999 8619
rect 15393 8585 15427 8619
rect 3617 8517 3651 8551
rect 5641 8517 5675 8551
rect 6101 8517 6135 8551
rect 9229 8517 9263 8551
rect 12265 8517 12299 8551
rect 15025 8517 15059 8551
rect 9459 8483 9493 8517
rect 2145 8449 2179 8483
rect 2329 8449 2363 8483
rect 2513 8449 2547 8483
rect 3341 8449 3375 8483
rect 3433 8449 3467 8483
rect 3709 8449 3743 8483
rect 3893 8449 3927 8483
rect 5365 8449 5399 8483
rect 5733 8449 5767 8483
rect 5917 8449 5951 8483
rect 6009 8449 6043 8483
rect 6193 8449 6227 8483
rect 7573 8449 7607 8483
rect 7941 8449 7975 8483
rect 8309 8449 8343 8483
rect 10057 8449 10091 8483
rect 10149 8449 10183 8483
rect 10425 8449 10459 8483
rect 11529 8449 11563 8483
rect 11713 8449 11747 8483
rect 11897 8449 11931 8483
rect 12081 8449 12115 8483
rect 14933 8449 14967 8483
rect 15209 8449 15243 8483
rect 1869 8381 1903 8415
rect 9689 8381 9723 8415
rect 10333 8381 10367 8415
rect 2789 8313 2823 8347
rect 3617 8313 3651 8347
rect 5641 8313 5675 8347
rect 8125 8313 8159 8347
rect 9597 8313 9631 8347
rect 10793 8313 10827 8347
rect 1961 8245 1995 8279
rect 3801 8245 3835 8279
rect 9413 8245 9447 8279
rect 12449 8245 12483 8279
rect 1685 8041 1719 8075
rect 2513 8041 2547 8075
rect 4629 8041 4663 8075
rect 8401 8041 8435 8075
rect 8585 8041 8619 8075
rect 12357 8041 12391 8075
rect 14749 8041 14783 8075
rect 5089 7973 5123 8007
rect 6929 7973 6963 8007
rect 13737 7973 13771 8007
rect 3157 7905 3191 7939
rect 9045 7905 9079 7939
rect 9689 7905 9723 7939
rect 12817 7905 12851 7939
rect 13277 7905 13311 7939
rect 14381 7905 14415 7939
rect 15209 7905 15243 7939
rect 15669 7905 15703 7939
rect 1777 7837 1811 7871
rect 1869 7837 1903 7871
rect 2237 7837 2271 7871
rect 2329 7837 2363 7871
rect 2697 7837 2731 7871
rect 3249 7837 3283 7871
rect 3801 7837 3835 7871
rect 4905 7837 4939 7871
rect 6837 7837 6871 7871
rect 6929 7837 6963 7871
rect 7113 7837 7147 7871
rect 7481 7837 7515 7871
rect 8309 7837 8343 7871
rect 8953 7837 8987 7871
rect 9229 7837 9263 7871
rect 9781 7837 9815 7871
rect 12081 7837 12115 7871
rect 12357 7837 12391 7871
rect 12725 7837 12759 7871
rect 12909 7837 12943 7871
rect 13369 7837 13403 7871
rect 14473 7837 14507 7871
rect 15301 7837 15335 7871
rect 15761 7837 15795 7871
rect 2027 7769 2061 7803
rect 2145 7769 2179 7803
rect 4597 7769 4631 7803
rect 4813 7769 4847 7803
rect 7297 7769 7331 7803
rect 7389 7769 7423 7803
rect 8769 7769 8803 7803
rect 9873 7769 9907 7803
rect 2881 7701 2915 7735
rect 3985 7701 4019 7735
rect 4445 7701 4479 7735
rect 7665 7701 7699 7735
rect 8125 7701 8159 7735
rect 8569 7701 8603 7735
rect 12173 7701 12207 7735
rect 15945 7701 15979 7735
rect 2329 7497 2363 7531
rect 2421 7497 2455 7531
rect 3709 7497 3743 7531
rect 4537 7497 4571 7531
rect 6101 7497 6135 7531
rect 9873 7497 9907 7531
rect 12465 7497 12499 7531
rect 12633 7497 12667 7531
rect 13645 7497 13679 7531
rect 14933 7497 14967 7531
rect 1501 7429 1535 7463
rect 1961 7429 1995 7463
rect 2881 7429 2915 7463
rect 3097 7429 3131 7463
rect 5641 7429 5675 7463
rect 5733 7429 5767 7463
rect 7481 7429 7515 7463
rect 8861 7429 8895 7463
rect 9505 7429 9539 7463
rect 9705 7429 9739 7463
rect 10333 7429 10367 7463
rect 11161 7429 11195 7463
rect 11345 7429 11379 7463
rect 12265 7429 12299 7463
rect 14473 7429 14507 7463
rect 1777 7361 1811 7395
rect 2053 7361 2087 7395
rect 2145 7361 2179 7395
rect 2421 7361 2455 7395
rect 2605 7361 2639 7395
rect 3901 7361 3935 7395
rect 4169 7361 4203 7395
rect 4445 7361 4479 7395
rect 4629 7361 4663 7395
rect 4721 7361 4755 7395
rect 4905 7361 4939 7395
rect 5549 7361 5583 7395
rect 5917 7361 5951 7395
rect 6009 7361 6043 7395
rect 6377 7361 6411 7395
rect 7297 7361 7331 7395
rect 7573 7361 7607 7395
rect 7670 7383 7704 7417
rect 9045 7361 9079 7395
rect 10149 7361 10183 7395
rect 10977 7361 11011 7395
rect 13185 7361 13219 7395
rect 1685 7293 1719 7327
rect 3985 7293 4019 7327
rect 7389 7293 7423 7327
rect 9229 7293 9263 7327
rect 3249 7225 3283 7259
rect 13461 7225 13495 7259
rect 14749 7225 14783 7259
rect 3065 7157 3099 7191
rect 4353 7157 4387 7191
rect 4813 7157 4847 7191
rect 5365 7157 5399 7191
rect 6561 7157 6595 7191
rect 9689 7157 9723 7191
rect 10517 7157 10551 7191
rect 12449 7157 12483 7191
rect 6101 6953 6135 6987
rect 9321 6953 9355 6987
rect 12173 6953 12207 6987
rect 3065 6885 3099 6919
rect 1777 6817 1811 6851
rect 6909 6817 6943 6851
rect 8033 6817 8067 6851
rect 2237 6749 2271 6783
rect 2973 6749 3007 6783
rect 3148 6749 3182 6783
rect 3249 6749 3283 6783
rect 4169 6749 4203 6783
rect 4537 6749 4571 6783
rect 4629 6749 4663 6783
rect 4997 6749 5031 6783
rect 5181 6749 5215 6783
rect 5457 6749 5491 6783
rect 5549 6749 5583 6783
rect 5825 6749 5859 6783
rect 5917 6749 5951 6783
rect 7113 6749 7147 6783
rect 7941 6749 7975 6783
rect 8125 6749 8159 6783
rect 8217 6749 8251 6783
rect 9505 6749 9539 6783
rect 9597 6749 9631 6783
rect 10701 6749 10735 6783
rect 10885 6749 10919 6783
rect 11805 6749 11839 6783
rect 11897 6749 11931 6783
rect 12081 6749 12115 6783
rect 12265 6749 12299 6783
rect 2513 6681 2547 6715
rect 5641 6681 5675 6715
rect 6837 6681 6871 6715
rect 9321 6681 9355 6715
rect 2789 6613 2823 6647
rect 3341 6613 3375 6647
rect 5089 6613 5123 6647
rect 5273 6613 5307 6647
rect 7021 6613 7055 6647
rect 8309 6613 8343 6647
rect 11713 6613 11747 6647
rect 2421 6409 2455 6443
rect 5549 6409 5583 6443
rect 7481 6409 7515 6443
rect 8217 6409 8251 6443
rect 8651 6409 8685 6443
rect 9045 6409 9079 6443
rect 12817 6409 12851 6443
rect 14841 6409 14875 6443
rect 3433 6341 3467 6375
rect 4629 6341 4663 6375
rect 4813 6341 4847 6375
rect 5029 6341 5063 6375
rect 8861 6341 8895 6375
rect 14473 6341 14507 6375
rect 1409 6273 1443 6307
rect 2237 6273 2271 6307
rect 2329 6273 2363 6307
rect 2881 6273 2915 6307
rect 3709 6273 3743 6307
rect 4445 6273 4479 6307
rect 5733 6273 5767 6307
rect 5917 6273 5951 6307
rect 6009 6273 6043 6307
rect 6377 6273 6411 6307
rect 6561 6273 6595 6307
rect 6653 6273 6687 6307
rect 6745 6273 6779 6307
rect 7849 6273 7883 6307
rect 8033 6273 8067 6307
rect 9229 6273 9263 6307
rect 11713 6273 11747 6307
rect 12817 6273 12851 6307
rect 13921 6273 13955 6307
rect 14105 6273 14139 6307
rect 14381 6273 14415 6307
rect 14657 6273 14691 6307
rect 1685 6205 1719 6239
rect 2605 6205 2639 6239
rect 2697 6205 2731 6239
rect 3893 6205 3927 6239
rect 7021 6205 7055 6239
rect 11621 6205 11655 6239
rect 12449 6205 12483 6239
rect 13001 6205 13035 6239
rect 14289 6205 14323 6239
rect 6929 6137 6963 6171
rect 1961 6069 1995 6103
rect 4261 6069 4295 6103
rect 4997 6069 5031 6103
rect 5181 6069 5215 6103
rect 7665 6069 7699 6103
rect 8493 6069 8527 6103
rect 8677 6069 8711 6103
rect 11989 6069 12023 6103
rect 3525 5865 3559 5899
rect 4813 5865 4847 5899
rect 6745 5865 6779 5899
rect 6929 5865 6963 5899
rect 7573 5865 7607 5899
rect 9137 5865 9171 5899
rect 11069 5865 11103 5899
rect 12633 5865 12667 5899
rect 14657 5865 14691 5899
rect 9321 5797 9355 5831
rect 9965 5797 9999 5831
rect 10609 5797 10643 5831
rect 11621 5797 11655 5831
rect 12127 5797 12161 5831
rect 2605 5729 2639 5763
rect 5917 5729 5951 5763
rect 7205 5729 7239 5763
rect 9505 5729 9539 5763
rect 10701 5729 10735 5763
rect 12357 5729 12391 5763
rect 13829 5729 13863 5763
rect 14197 5729 14231 5763
rect 14841 5729 14875 5763
rect 15301 5729 15335 5763
rect 1593 5661 1627 5695
rect 1869 5661 1903 5695
rect 1961 5661 1995 5695
rect 2237 5661 2271 5695
rect 2513 5661 2547 5695
rect 2789 5661 2823 5695
rect 3065 5661 3099 5695
rect 3341 5661 3375 5695
rect 3893 5661 3927 5695
rect 4077 5661 4111 5695
rect 4540 5661 4574 5695
rect 4813 5661 4847 5695
rect 6009 5661 6043 5695
rect 6101 5661 6135 5695
rect 6193 5661 6227 5695
rect 7113 5661 7147 5695
rect 7297 5661 7331 5695
rect 7389 5661 7423 5695
rect 8033 5661 8067 5695
rect 9597 5661 9631 5695
rect 10425 5661 10459 5695
rect 10609 5661 10643 5695
rect 10885 5661 10919 5695
rect 11437 5661 11471 5695
rect 11529 5661 11563 5695
rect 11713 5661 11747 5695
rect 12219 5661 12253 5695
rect 13093 5661 13127 5695
rect 13369 5661 13403 5695
rect 14289 5661 14323 5695
rect 14933 5661 14967 5695
rect 15669 5661 15703 5695
rect 1777 5593 1811 5627
rect 3985 5593 4019 5627
rect 4629 5593 4663 5627
rect 6561 5593 6595 5627
rect 6761 5593 6795 5627
rect 8953 5593 8987 5627
rect 9153 5593 9187 5627
rect 11989 5593 12023 5627
rect 2145 5525 2179 5559
rect 6377 5525 6411 5559
rect 8217 5525 8251 5559
rect 11897 5525 11931 5559
rect 15945 5525 15979 5559
rect 13277 5321 13311 5355
rect 2421 5253 2455 5287
rect 2697 5253 2731 5287
rect 2881 5253 2915 5287
rect 7849 5253 7883 5287
rect 7941 5253 7975 5287
rect 11529 5253 11563 5287
rect 11713 5253 11747 5287
rect 1869 5185 1903 5219
rect 4169 5185 4203 5219
rect 4261 5185 4295 5219
rect 4445 5185 4479 5219
rect 6377 5185 6411 5219
rect 6653 5185 6687 5219
rect 7481 5185 7515 5219
rect 7665 5185 7699 5219
rect 8033 5185 8067 5219
rect 8493 5185 8527 5219
rect 8585 5185 8619 5219
rect 8769 5185 8803 5219
rect 9137 5185 9171 5219
rect 9229 5185 9263 5219
rect 9406 5185 9440 5219
rect 9965 5185 9999 5219
rect 10793 5185 10827 5219
rect 12817 5185 12851 5219
rect 13185 5185 13219 5219
rect 3801 5117 3835 5151
rect 5365 5117 5399 5151
rect 8861 5117 8895 5151
rect 8217 5049 8251 5083
rect 9045 5049 9079 5083
rect 9321 5049 9355 5083
rect 3985 4981 4019 5015
rect 7297 4981 7331 5015
rect 8769 4981 8803 5015
rect 8953 4981 8987 5015
rect 10057 4981 10091 5015
rect 10425 4981 10459 5015
rect 10609 4981 10643 5015
rect 11897 4981 11931 5015
rect 2973 4777 3007 4811
rect 6009 4777 6043 4811
rect 11437 4777 11471 4811
rect 6285 4709 6319 4743
rect 11253 4709 11287 4743
rect 1777 4641 1811 4675
rect 2697 4641 2731 4675
rect 5825 4641 5859 4675
rect 7481 4641 7515 4675
rect 8309 4641 8343 4675
rect 10425 4641 10459 4675
rect 10885 4641 10919 4675
rect 1501 4573 1535 4607
rect 2237 4573 2271 4607
rect 2513 4573 2547 4607
rect 3249 4573 3283 4607
rect 3433 4573 3467 4607
rect 3525 4573 3559 4607
rect 4169 4573 4203 4607
rect 6101 4573 6135 4607
rect 6193 4573 6227 4607
rect 6469 4573 6503 4607
rect 7389 4573 7423 4607
rect 7757 4573 7791 4607
rect 7849 4573 7883 4607
rect 10517 4573 10551 4607
rect 2329 4505 2363 4539
rect 2789 4505 2823 4539
rect 2989 4505 3023 4539
rect 6929 4505 6963 4539
rect 7021 4505 7055 4539
rect 10977 4505 11011 4539
rect 3157 4437 3191 4471
rect 3341 4437 3375 4471
rect 4353 4437 4387 4471
rect 5825 4437 5859 4471
rect 7665 4437 7699 4471
rect 2145 4233 2179 4267
rect 3617 4233 3651 4267
rect 2053 4165 2087 4199
rect 2789 4165 2823 4199
rect 2881 4165 2915 4199
rect 3249 4165 3283 4199
rect 3433 4165 3467 4199
rect 1409 4097 1443 4131
rect 1685 4097 1719 4131
rect 2605 4097 2639 4131
rect 2973 4097 3007 4131
rect 3525 4097 3559 4131
rect 4169 4097 4203 4131
rect 7389 4097 7423 4131
rect 8769 4097 8803 4131
rect 9229 4097 9263 4131
rect 11529 4097 11563 4131
rect 11713 4097 11747 4131
rect 11989 4097 12023 4131
rect 12449 4097 12483 4131
rect 12541 4097 12575 4131
rect 12725 4097 12759 4131
rect 12909 4097 12943 4131
rect 13737 4097 13771 4131
rect 14013 4097 14047 4131
rect 14105 4097 14139 4131
rect 14289 4097 14323 4131
rect 14473 4097 14507 4131
rect 4261 4029 4295 4063
rect 7481 4029 7515 4063
rect 7757 4029 7791 4063
rect 8677 4029 8711 4063
rect 12081 4029 12115 4063
rect 13553 4029 13587 4063
rect 13921 4029 13955 4063
rect 11529 3961 11563 3995
rect 3157 3893 3191 3927
rect 3801 3893 3835 3927
rect 4445 3893 4479 3927
rect 9137 3893 9171 3927
rect 9321 3893 9355 3927
rect 9689 3893 9723 3927
rect 12357 3893 12391 3927
rect 6377 3689 6411 3723
rect 9413 3689 9447 3723
rect 13921 3689 13955 3723
rect 6745 3621 6779 3655
rect 15945 3621 15979 3655
rect 1685 3553 1719 3587
rect 9597 3553 9631 3587
rect 12633 3553 12667 3587
rect 13093 3553 13127 3587
rect 13645 3553 13679 3587
rect 14197 3553 14231 3587
rect 14657 3553 14691 3587
rect 1409 3485 1443 3519
rect 4353 3485 4387 3519
rect 5825 3485 5859 3519
rect 5917 3485 5951 3519
rect 6193 3485 6227 3519
rect 6469 3485 6503 3519
rect 6653 3485 6687 3519
rect 6745 3485 6779 3519
rect 6929 3485 6963 3519
rect 8125 3485 8159 3519
rect 9321 3485 9355 3519
rect 12725 3485 12759 3519
rect 13553 3485 13587 3519
rect 14289 3485 14323 3519
rect 15761 3485 15795 3519
rect 6561 3417 6595 3451
rect 9597 3417 9631 3451
rect 4169 3349 4203 3383
rect 5641 3349 5675 3383
rect 6009 3349 6043 3383
rect 7941 3349 7975 3383
rect 4261 3145 4295 3179
rect 6193 3145 6227 3179
rect 7021 3145 7055 3179
rect 8325 3145 8359 3179
rect 12081 3145 12115 3179
rect 7205 3077 7239 3111
rect 7389 3077 7423 3111
rect 7665 3077 7699 3111
rect 7865 3077 7899 3111
rect 8125 3077 8159 3111
rect 1409 3009 1443 3043
rect 2973 3009 3007 3043
rect 3709 3009 3743 3043
rect 4169 3009 4203 3043
rect 4445 3009 4479 3043
rect 5181 3009 5215 3043
rect 5825 3009 5859 3043
rect 6929 3009 6963 3043
rect 7297 3009 7331 3043
rect 7573 3009 7607 3043
rect 8585 3009 8619 3043
rect 8769 3009 8803 3043
rect 8861 3009 8895 3043
rect 8953 3009 8987 3043
rect 9413 3009 9447 3043
rect 10241 3009 10275 3043
rect 11161 3009 11195 3043
rect 11345 3009 11379 3043
rect 11713 3009 11747 3043
rect 12173 3009 12207 3043
rect 1961 2941 1995 2975
rect 3433 2941 3467 2975
rect 3617 2941 3651 2975
rect 5273 2941 5307 2975
rect 5733 2941 5767 2975
rect 9321 2941 9355 2975
rect 10333 2941 10367 2975
rect 11621 2941 11655 2975
rect 4077 2873 4111 2907
rect 5549 2873 5583 2907
rect 7573 2873 7607 2907
rect 8033 2873 8067 2907
rect 9781 2873 9815 2907
rect 10609 2873 10643 2907
rect 12265 2873 12299 2907
rect 3249 2805 3283 2839
rect 4629 2805 4663 2839
rect 7205 2805 7239 2839
rect 7849 2805 7883 2839
rect 8309 2805 8343 2839
rect 8493 2805 8527 2839
rect 8585 2805 8619 2839
rect 10885 2805 10919 2839
rect 11161 2805 11195 2839
rect 7389 2601 7423 2635
rect 7757 2601 7791 2635
rect 8033 2601 8067 2635
rect 9321 2601 9355 2635
rect 10517 2601 10551 2635
rect 4721 2397 4755 2431
rect 7205 2397 7239 2431
rect 7757 2397 7791 2431
rect 7941 2397 7975 2431
rect 8217 2397 8251 2431
rect 8677 2397 8711 2431
rect 9137 2397 9171 2431
rect 10333 2397 10367 2431
rect 10517 2397 10551 2431
rect 12449 2397 12483 2431
rect 4813 2261 4847 2295
rect 8401 2261 8435 2295
rect 12541 2261 12575 2295
<< metal1 >>
rect 1104 17434 16376 17456
rect 1104 17382 3519 17434
rect 3571 17382 3583 17434
rect 3635 17382 3647 17434
rect 3699 17382 3711 17434
rect 3763 17382 3775 17434
rect 3827 17382 7337 17434
rect 7389 17382 7401 17434
rect 7453 17382 7465 17434
rect 7517 17382 7529 17434
rect 7581 17382 7593 17434
rect 7645 17382 11155 17434
rect 11207 17382 11219 17434
rect 11271 17382 11283 17434
rect 11335 17382 11347 17434
rect 11399 17382 11411 17434
rect 11463 17382 14973 17434
rect 15025 17382 15037 17434
rect 15089 17382 15101 17434
rect 15153 17382 15165 17434
rect 15217 17382 15229 17434
rect 15281 17382 16376 17434
rect 1104 17360 16376 17382
rect 13814 17280 13820 17332
rect 13872 17320 13878 17332
rect 14277 17323 14335 17329
rect 14277 17320 14289 17323
rect 13872 17292 14289 17320
rect 13872 17280 13878 17292
rect 14277 17289 14289 17292
rect 14323 17289 14335 17323
rect 14277 17283 14335 17289
rect 14826 17280 14832 17332
rect 14884 17320 14890 17332
rect 15289 17323 15347 17329
rect 15289 17320 15301 17323
rect 14884 17292 15301 17320
rect 14884 17280 14890 17292
rect 15289 17289 15301 17292
rect 15335 17289 15347 17323
rect 15289 17283 15347 17289
rect 12434 17212 12440 17264
rect 12492 17252 12498 17264
rect 12529 17255 12587 17261
rect 12529 17252 12541 17255
rect 12492 17224 12541 17252
rect 12492 17212 12498 17224
rect 12529 17221 12541 17224
rect 12575 17221 12587 17255
rect 12529 17215 12587 17221
rect 7190 17144 7196 17196
rect 7248 17144 7254 17196
rect 7282 17144 7288 17196
rect 7340 17184 7346 17196
rect 7377 17187 7435 17193
rect 7377 17184 7389 17187
rect 7340 17156 7389 17184
rect 7340 17144 7346 17156
rect 7377 17153 7389 17156
rect 7423 17184 7435 17187
rect 8018 17184 8024 17196
rect 7423 17156 8024 17184
rect 7423 17153 7435 17156
rect 7377 17147 7435 17153
rect 8018 17144 8024 17156
rect 8076 17144 8082 17196
rect 10318 17144 10324 17196
rect 10376 17144 10382 17196
rect 10410 17144 10416 17196
rect 10468 17144 10474 17196
rect 10597 17187 10655 17193
rect 10597 17153 10609 17187
rect 10643 17153 10655 17187
rect 10597 17147 10655 17153
rect 9858 17076 9864 17128
rect 9916 17116 9922 17128
rect 10612 17116 10640 17147
rect 12158 17144 12164 17196
rect 12216 17144 12222 17196
rect 12802 17144 12808 17196
rect 12860 17184 12866 17196
rect 12897 17187 12955 17193
rect 12897 17184 12909 17187
rect 12860 17156 12909 17184
rect 12860 17144 12866 17156
rect 12897 17153 12909 17156
rect 12943 17153 12955 17187
rect 12897 17147 12955 17153
rect 13081 17187 13139 17193
rect 13081 17153 13093 17187
rect 13127 17153 13139 17187
rect 13081 17147 13139 17153
rect 10870 17116 10876 17128
rect 9916 17088 10876 17116
rect 9916 17076 9922 17088
rect 10870 17076 10876 17088
rect 10928 17076 10934 17128
rect 12066 17076 12072 17128
rect 12124 17116 12130 17128
rect 13096 17116 13124 17147
rect 14182 17144 14188 17196
rect 14240 17144 14246 17196
rect 15010 17144 15016 17196
rect 15068 17144 15074 17196
rect 12124 17088 13124 17116
rect 12124 17076 12130 17088
rect 7466 17008 7472 17060
rect 7524 17048 7530 17060
rect 12618 17048 12624 17060
rect 7524 17020 12624 17048
rect 7524 17008 7530 17020
rect 12618 17008 12624 17020
rect 12676 17008 12682 17060
rect 7561 16983 7619 16989
rect 7561 16949 7573 16983
rect 7607 16980 7619 16983
rect 9030 16980 9036 16992
rect 7607 16952 9036 16980
rect 7607 16949 7619 16952
rect 7561 16943 7619 16949
rect 9030 16940 9036 16952
rect 9088 16940 9094 16992
rect 10597 16983 10655 16989
rect 10597 16949 10609 16983
rect 10643 16980 10655 16983
rect 11606 16980 11612 16992
rect 10643 16952 11612 16980
rect 10643 16949 10655 16952
rect 10597 16943 10655 16949
rect 11606 16940 11612 16952
rect 11664 16940 11670 16992
rect 12894 16940 12900 16992
rect 12952 16940 12958 16992
rect 1104 16890 16376 16912
rect 1104 16838 2859 16890
rect 2911 16838 2923 16890
rect 2975 16838 2987 16890
rect 3039 16838 3051 16890
rect 3103 16838 3115 16890
rect 3167 16838 6677 16890
rect 6729 16838 6741 16890
rect 6793 16838 6805 16890
rect 6857 16838 6869 16890
rect 6921 16838 6933 16890
rect 6985 16838 10495 16890
rect 10547 16838 10559 16890
rect 10611 16838 10623 16890
rect 10675 16838 10687 16890
rect 10739 16838 10751 16890
rect 10803 16838 14313 16890
rect 14365 16838 14377 16890
rect 14429 16838 14441 16890
rect 14493 16838 14505 16890
rect 14557 16838 14569 16890
rect 14621 16838 16376 16890
rect 1104 16816 16376 16838
rect 6641 16779 6699 16785
rect 6641 16745 6653 16779
rect 6687 16776 6699 16779
rect 7190 16776 7196 16788
rect 6687 16748 7196 16776
rect 6687 16745 6699 16748
rect 6641 16739 6699 16745
rect 7190 16736 7196 16748
rect 7248 16736 7254 16788
rect 7466 16736 7472 16788
rect 7524 16736 7530 16788
rect 8018 16736 8024 16788
rect 8076 16776 8082 16788
rect 8076 16748 8524 16776
rect 8076 16736 8082 16748
rect 5994 16532 6000 16584
rect 6052 16572 6058 16584
rect 6365 16575 6423 16581
rect 6365 16572 6377 16575
rect 6052 16544 6377 16572
rect 6052 16532 6058 16544
rect 6365 16541 6377 16544
rect 6411 16572 6423 16575
rect 6917 16575 6975 16581
rect 6917 16572 6929 16575
rect 6411 16544 6929 16572
rect 6411 16541 6423 16544
rect 6365 16535 6423 16541
rect 6917 16541 6929 16544
rect 6963 16541 6975 16575
rect 6917 16535 6975 16541
rect 7190 16532 7196 16584
rect 7248 16572 7254 16584
rect 7285 16575 7343 16581
rect 7285 16572 7297 16575
rect 7248 16544 7297 16572
rect 7248 16532 7254 16544
rect 7285 16541 7297 16544
rect 7331 16541 7343 16575
rect 7285 16535 7343 16541
rect 7377 16575 7435 16581
rect 7377 16541 7389 16575
rect 7423 16541 7435 16575
rect 7484 16572 7512 16736
rect 8297 16711 8355 16717
rect 8297 16708 8309 16711
rect 7760 16680 8309 16708
rect 7760 16581 7788 16680
rect 8297 16677 8309 16680
rect 8343 16677 8355 16711
rect 8297 16671 8355 16677
rect 8202 16640 8208 16652
rect 7852 16612 8208 16640
rect 7852 16581 7880 16612
rect 8202 16600 8208 16612
rect 8260 16600 8266 16652
rect 7561 16575 7619 16581
rect 7561 16572 7573 16575
rect 7484 16544 7573 16572
rect 7377 16535 7435 16541
rect 7561 16541 7573 16544
rect 7607 16541 7619 16575
rect 7561 16535 7619 16541
rect 7745 16575 7803 16581
rect 7745 16541 7757 16575
rect 7791 16541 7803 16575
rect 7745 16535 7803 16541
rect 7837 16575 7895 16581
rect 7837 16541 7849 16575
rect 7883 16541 7895 16575
rect 7837 16535 7895 16541
rect 6546 16464 6552 16516
rect 6604 16504 6610 16516
rect 6641 16507 6699 16513
rect 6641 16504 6653 16507
rect 6604 16476 6653 16504
rect 6604 16464 6610 16476
rect 6641 16473 6653 16476
rect 6687 16473 6699 16507
rect 7392 16504 7420 16535
rect 7926 16532 7932 16584
rect 7984 16532 7990 16584
rect 8018 16532 8024 16584
rect 8076 16532 8082 16584
rect 8496 16581 8524 16748
rect 9030 16736 9036 16788
rect 9088 16776 9094 16788
rect 9677 16779 9735 16785
rect 9677 16776 9689 16779
rect 9088 16748 9689 16776
rect 9088 16736 9094 16748
rect 9677 16745 9689 16748
rect 9723 16745 9735 16779
rect 9677 16739 9735 16745
rect 10134 16736 10140 16788
rect 10192 16776 10198 16788
rect 10229 16779 10287 16785
rect 10229 16776 10241 16779
rect 10192 16748 10241 16776
rect 10192 16736 10198 16748
rect 10229 16745 10241 16748
rect 10275 16745 10287 16779
rect 10229 16739 10287 16745
rect 10410 16736 10416 16788
rect 10468 16736 10474 16788
rect 10502 16736 10508 16788
rect 10560 16776 10566 16788
rect 10873 16779 10931 16785
rect 10873 16776 10885 16779
rect 10560 16748 10885 16776
rect 10560 16736 10566 16748
rect 10873 16745 10885 16748
rect 10919 16745 10931 16779
rect 10873 16739 10931 16745
rect 11885 16779 11943 16785
rect 11885 16745 11897 16779
rect 11931 16745 11943 16779
rect 11885 16739 11943 16745
rect 9048 16649 9076 16736
rect 9493 16711 9551 16717
rect 9493 16677 9505 16711
rect 9539 16677 9551 16711
rect 9493 16671 9551 16677
rect 10045 16711 10103 16717
rect 10045 16677 10057 16711
rect 10091 16708 10103 16711
rect 10428 16708 10456 16736
rect 10091 16680 10456 16708
rect 10091 16677 10103 16680
rect 10045 16671 10103 16677
rect 9033 16643 9091 16649
rect 9033 16609 9045 16643
rect 9079 16609 9091 16643
rect 9508 16640 9536 16671
rect 9508 16612 10272 16640
rect 9033 16603 9091 16609
rect 10244 16584 10272 16612
rect 8297 16575 8355 16581
rect 8297 16572 8309 16575
rect 8128 16544 8309 16572
rect 8128 16504 8156 16544
rect 8297 16541 8309 16544
rect 8343 16541 8355 16575
rect 8297 16535 8355 16541
rect 8481 16575 8539 16581
rect 8481 16541 8493 16575
rect 8527 16541 8539 16575
rect 8481 16535 8539 16541
rect 8938 16532 8944 16584
rect 8996 16572 9002 16584
rect 9125 16575 9183 16581
rect 9125 16572 9137 16575
rect 8996 16544 9137 16572
rect 8996 16532 9002 16544
rect 9125 16541 9137 16544
rect 9171 16572 9183 16575
rect 9585 16575 9643 16581
rect 9585 16572 9597 16575
rect 9171 16544 9597 16572
rect 9171 16541 9183 16544
rect 9125 16535 9183 16541
rect 9585 16541 9597 16544
rect 9631 16541 9643 16575
rect 9585 16535 9643 16541
rect 10226 16532 10232 16584
rect 10284 16532 10290 16584
rect 10318 16532 10324 16584
rect 10376 16532 10382 16584
rect 7392 16476 8156 16504
rect 10428 16504 10456 16680
rect 10888 16640 10916 16739
rect 11517 16711 11575 16717
rect 11517 16677 11529 16711
rect 11563 16708 11575 16711
rect 11900 16708 11928 16739
rect 12066 16736 12072 16788
rect 12124 16736 12130 16788
rect 12158 16736 12164 16788
rect 12216 16736 12222 16788
rect 13357 16779 13415 16785
rect 13357 16745 13369 16779
rect 13403 16776 13415 16779
rect 14182 16776 14188 16788
rect 13403 16748 14188 16776
rect 13403 16745 13415 16748
rect 13357 16739 13415 16745
rect 14182 16736 14188 16748
rect 14240 16736 14246 16788
rect 14553 16779 14611 16785
rect 14553 16745 14565 16779
rect 14599 16776 14611 16779
rect 15010 16776 15016 16788
rect 14599 16748 15016 16776
rect 14599 16745 14611 16748
rect 14553 16739 14611 16745
rect 15010 16736 15016 16748
rect 15068 16736 15074 16788
rect 12526 16708 12532 16720
rect 11563 16680 12532 16708
rect 11563 16677 11575 16680
rect 11517 16671 11575 16677
rect 12526 16668 12532 16680
rect 12584 16668 12590 16720
rect 11149 16643 11207 16649
rect 11149 16640 11161 16643
rect 10888 16612 11161 16640
rect 11149 16609 11161 16612
rect 11195 16609 11207 16643
rect 12894 16640 12900 16652
rect 11149 16603 11207 16609
rect 12452 16612 12900 16640
rect 12359 16585 12417 16591
rect 11333 16575 11391 16581
rect 11333 16572 11345 16575
rect 10796 16544 11345 16572
rect 10689 16507 10747 16513
rect 10689 16504 10701 16507
rect 10428 16476 10701 16504
rect 6641 16467 6699 16473
rect 7760 16448 7788 16476
rect 10689 16473 10701 16476
rect 10735 16473 10747 16507
rect 10689 16467 10747 16473
rect 6454 16396 6460 16448
rect 6512 16396 6518 16448
rect 7742 16396 7748 16448
rect 7800 16396 7806 16448
rect 8205 16439 8263 16445
rect 8205 16405 8217 16439
rect 8251 16436 8263 16439
rect 9858 16436 9864 16448
rect 8251 16408 9864 16436
rect 8251 16405 8263 16408
rect 8205 16399 8263 16405
rect 9858 16396 9864 16408
rect 9916 16396 9922 16448
rect 10597 16439 10655 16445
rect 10597 16405 10609 16439
rect 10643 16436 10655 16439
rect 10796 16436 10824 16544
rect 11333 16541 11345 16544
rect 11379 16541 11391 16575
rect 12359 16551 12371 16585
rect 12405 16582 12417 16585
rect 12452 16582 12480 16612
rect 12894 16600 12900 16612
rect 12952 16600 12958 16652
rect 14366 16600 14372 16652
rect 14424 16600 14430 16652
rect 12405 16554 12480 16582
rect 12510 16575 12568 16581
rect 12405 16551 12417 16554
rect 12359 16545 12417 16551
rect 11333 16535 11391 16541
rect 12510 16541 12522 16575
rect 12556 16572 12568 16575
rect 12556 16541 12572 16572
rect 12510 16535 12572 16541
rect 10870 16464 10876 16516
rect 10928 16513 10934 16516
rect 10928 16507 10947 16513
rect 10935 16473 10947 16507
rect 10928 16467 10947 16473
rect 11701 16507 11759 16513
rect 11701 16473 11713 16507
rect 11747 16504 11759 16507
rect 12544 16504 12572 16535
rect 12618 16532 12624 16584
rect 12676 16532 12682 16584
rect 12710 16532 12716 16584
rect 12768 16532 12774 16584
rect 12989 16575 13047 16581
rect 12989 16541 13001 16575
rect 13035 16572 13047 16575
rect 13035 16544 13676 16572
rect 13035 16541 13047 16544
rect 12989 16535 13047 16541
rect 13004 16504 13032 16535
rect 11747 16476 12434 16504
rect 12544 16476 13032 16504
rect 11747 16473 11759 16476
rect 11701 16467 11759 16473
rect 10928 16464 10934 16467
rect 10643 16408 10824 16436
rect 10643 16405 10655 16408
rect 10597 16399 10655 16405
rect 11054 16396 11060 16448
rect 11112 16396 11118 16448
rect 11882 16396 11888 16448
rect 11940 16445 11946 16448
rect 11940 16439 11959 16445
rect 11947 16405 11959 16439
rect 12406 16436 12434 16476
rect 13648 16448 13676 16544
rect 13722 16532 13728 16584
rect 13780 16572 13786 16584
rect 14277 16575 14335 16581
rect 14277 16572 14289 16575
rect 13780 16544 14289 16572
rect 13780 16532 13786 16544
rect 14277 16541 14289 16544
rect 14323 16541 14335 16575
rect 14277 16535 14335 16541
rect 12894 16436 12900 16448
rect 12406 16408 12900 16436
rect 11940 16399 11959 16405
rect 11940 16396 11946 16399
rect 12894 16396 12900 16408
rect 12952 16396 12958 16448
rect 13630 16396 13636 16448
rect 13688 16396 13694 16448
rect 1104 16346 16376 16368
rect 1104 16294 3519 16346
rect 3571 16294 3583 16346
rect 3635 16294 3647 16346
rect 3699 16294 3711 16346
rect 3763 16294 3775 16346
rect 3827 16294 7337 16346
rect 7389 16294 7401 16346
rect 7453 16294 7465 16346
rect 7517 16294 7529 16346
rect 7581 16294 7593 16346
rect 7645 16294 11155 16346
rect 11207 16294 11219 16346
rect 11271 16294 11283 16346
rect 11335 16294 11347 16346
rect 11399 16294 11411 16346
rect 11463 16294 14973 16346
rect 15025 16294 15037 16346
rect 15089 16294 15101 16346
rect 15153 16294 15165 16346
rect 15217 16294 15229 16346
rect 15281 16294 16376 16346
rect 1104 16272 16376 16294
rect 5813 16235 5871 16241
rect 5813 16201 5825 16235
rect 5859 16232 5871 16235
rect 7653 16235 7711 16241
rect 5859 16204 7328 16232
rect 5859 16201 5871 16204
rect 5813 16195 5871 16201
rect 7300 16173 7328 16204
rect 7653 16201 7665 16235
rect 7699 16232 7711 16235
rect 7742 16232 7748 16244
rect 7699 16204 7748 16232
rect 7699 16201 7711 16204
rect 7653 16195 7711 16201
rect 7742 16192 7748 16204
rect 7800 16192 7806 16244
rect 11609 16235 11667 16241
rect 11609 16201 11621 16235
rect 11655 16232 11667 16235
rect 11882 16232 11888 16244
rect 11655 16204 11888 16232
rect 11655 16201 11667 16204
rect 11609 16195 11667 16201
rect 11882 16192 11888 16204
rect 11940 16232 11946 16244
rect 12529 16235 12587 16241
rect 11940 16204 12434 16232
rect 11940 16192 11946 16204
rect 5721 16167 5779 16173
rect 5721 16164 5733 16167
rect 4172 16136 5733 16164
rect 4172 16108 4200 16136
rect 5721 16133 5733 16136
rect 5767 16133 5779 16167
rect 6641 16167 6699 16173
rect 6641 16164 6653 16167
rect 5721 16127 5779 16133
rect 6012 16136 6653 16164
rect 4154 16056 4160 16108
rect 4212 16056 4218 16108
rect 5626 16056 5632 16108
rect 5684 16056 5690 16108
rect 5736 16028 5764 16127
rect 6012 16105 6040 16136
rect 6641 16133 6653 16136
rect 6687 16164 6699 16167
rect 7285 16167 7343 16173
rect 6687 16136 7144 16164
rect 6687 16133 6699 16136
rect 6641 16127 6699 16133
rect 7116 16108 7144 16136
rect 7285 16133 7297 16167
rect 7331 16133 7343 16167
rect 7285 16127 7343 16133
rect 5997 16099 6055 16105
rect 6549 16102 6607 16105
rect 5997 16065 6009 16099
rect 6043 16065 6055 16099
rect 5997 16059 6055 16065
rect 6472 16099 6607 16102
rect 6472 16074 6561 16099
rect 6472 16028 6500 16074
rect 6549 16065 6561 16074
rect 6595 16065 6607 16099
rect 6549 16059 6607 16065
rect 6733 16099 6791 16105
rect 6733 16065 6745 16099
rect 6779 16096 6791 16099
rect 6822 16096 6828 16108
rect 6779 16068 6828 16096
rect 6779 16065 6791 16068
rect 6733 16059 6791 16065
rect 6822 16056 6828 16068
rect 6880 16056 6886 16108
rect 6917 16099 6975 16105
rect 6917 16065 6929 16099
rect 6963 16065 6975 16099
rect 6917 16059 6975 16065
rect 6932 16028 6960 16059
rect 7098 16056 7104 16108
rect 7156 16056 7162 16108
rect 7300 16096 7328 16127
rect 7466 16124 7472 16176
rect 7524 16173 7530 16176
rect 7524 16167 7543 16173
rect 7531 16133 7543 16167
rect 7524 16127 7543 16133
rect 7524 16124 7530 16127
rect 8202 16124 8208 16176
rect 8260 16124 8266 16176
rect 10318 16124 10324 16176
rect 10376 16124 10382 16176
rect 12066 16124 12072 16176
rect 12124 16164 12130 16176
rect 12161 16167 12219 16173
rect 12161 16164 12173 16167
rect 12124 16136 12173 16164
rect 12124 16124 12130 16136
rect 12161 16133 12173 16136
rect 12207 16133 12219 16167
rect 12406 16164 12434 16204
rect 12529 16201 12541 16235
rect 12575 16232 12587 16235
rect 12710 16232 12716 16244
rect 12575 16204 12716 16232
rect 12575 16201 12587 16204
rect 12529 16195 12587 16201
rect 12710 16192 12716 16204
rect 12768 16192 12774 16244
rect 12805 16235 12863 16241
rect 12805 16201 12817 16235
rect 12851 16232 12863 16235
rect 12894 16232 12900 16244
rect 12851 16204 12900 16232
rect 12851 16201 12863 16204
rect 12805 16195 12863 16201
rect 12894 16192 12900 16204
rect 12952 16192 12958 16244
rect 13630 16192 13636 16244
rect 13688 16192 13694 16244
rect 12621 16167 12679 16173
rect 12621 16164 12633 16167
rect 12406 16136 12633 16164
rect 12161 16127 12219 16133
rect 12621 16133 12633 16136
rect 12667 16133 12679 16167
rect 13722 16164 13728 16176
rect 12621 16127 12679 16133
rect 12912 16136 13728 16164
rect 8220 16096 8248 16124
rect 7300 16068 8248 16096
rect 10045 16099 10103 16105
rect 7300 16028 7328 16068
rect 10045 16065 10057 16099
rect 10091 16096 10103 16099
rect 10336 16096 10364 16124
rect 10091 16068 10364 16096
rect 10091 16065 10103 16068
rect 10045 16059 10103 16065
rect 11054 16056 11060 16108
rect 11112 16096 11118 16108
rect 11517 16099 11575 16105
rect 11517 16096 11529 16099
rect 11112 16068 11529 16096
rect 11112 16056 11118 16068
rect 11517 16065 11529 16068
rect 11563 16065 11575 16099
rect 11517 16059 11575 16065
rect 11606 16056 11612 16108
rect 11664 16096 11670 16108
rect 11701 16099 11759 16105
rect 11701 16096 11713 16099
rect 11664 16068 11713 16096
rect 11664 16056 11670 16068
rect 11701 16065 11713 16068
rect 11747 16096 11759 16099
rect 12345 16099 12403 16105
rect 12345 16096 12357 16099
rect 11747 16068 12357 16096
rect 11747 16065 11759 16068
rect 11701 16059 11759 16065
rect 12345 16065 12357 16068
rect 12391 16065 12403 16099
rect 12345 16059 12403 16065
rect 12526 16056 12532 16108
rect 12584 16056 12590 16108
rect 12912 16105 12940 16136
rect 13722 16124 13728 16136
rect 13780 16173 13786 16176
rect 13780 16167 13843 16173
rect 13780 16133 13797 16167
rect 13831 16133 13843 16167
rect 13780 16127 13843 16133
rect 13780 16124 13786 16127
rect 13906 16124 13912 16176
rect 13964 16164 13970 16176
rect 14001 16167 14059 16173
rect 14001 16164 14013 16167
rect 13964 16136 14013 16164
rect 13964 16124 13970 16136
rect 14001 16133 14013 16136
rect 14047 16164 14059 16167
rect 14185 16167 14243 16173
rect 14185 16164 14197 16167
rect 14047 16136 14197 16164
rect 14047 16133 14059 16136
rect 14001 16127 14059 16133
rect 14185 16133 14197 16136
rect 14231 16133 14243 16167
rect 14185 16127 14243 16133
rect 12897 16099 12955 16105
rect 12897 16065 12909 16099
rect 12943 16065 12955 16099
rect 14093 16099 14151 16105
rect 14093 16096 14105 16099
rect 12897 16059 12955 16065
rect 13832 16068 14105 16096
rect 5736 16000 6868 16028
rect 6932 16000 7328 16028
rect 5905 15963 5963 15969
rect 5905 15929 5917 15963
rect 5951 15960 5963 15963
rect 5994 15960 6000 15972
rect 5951 15932 6000 15960
rect 5951 15929 5963 15932
rect 5905 15923 5963 15929
rect 5994 15920 6000 15932
rect 6052 15920 6058 15972
rect 6365 15963 6423 15969
rect 6365 15929 6377 15963
rect 6411 15960 6423 15963
rect 6454 15960 6460 15972
rect 6411 15932 6460 15960
rect 6411 15929 6423 15932
rect 6365 15923 6423 15929
rect 6454 15920 6460 15932
rect 6512 15920 6518 15972
rect 6840 15892 6868 16000
rect 10226 15988 10232 16040
rect 10284 16028 10290 16040
rect 10321 16031 10379 16037
rect 10321 16028 10333 16031
rect 10284 16000 10333 16028
rect 10284 15988 10290 16000
rect 10321 15997 10333 16000
rect 10367 15997 10379 16031
rect 12544 16028 12572 16056
rect 12912 16028 12940 16059
rect 12544 16000 12940 16028
rect 10321 15991 10379 15997
rect 10134 15920 10140 15972
rect 10192 15920 10198 15972
rect 12621 15963 12679 15969
rect 12621 15929 12633 15963
rect 12667 15960 12679 15963
rect 12802 15960 12808 15972
rect 12667 15932 12808 15960
rect 12667 15929 12679 15932
rect 12621 15923 12679 15929
rect 12802 15920 12808 15932
rect 12860 15920 12866 15972
rect 13832 15904 13860 16068
rect 14093 16065 14105 16068
rect 14139 16065 14151 16099
rect 14369 16099 14427 16105
rect 14369 16096 14381 16099
rect 14093 16059 14151 16065
rect 14200 16068 14381 16096
rect 14200 15904 14228 16068
rect 14369 16065 14381 16068
rect 14415 16065 14427 16099
rect 14369 16059 14427 16065
rect 14366 15920 14372 15972
rect 14424 15920 14430 15972
rect 7469 15895 7527 15901
rect 7469 15892 7481 15895
rect 6840 15864 7481 15892
rect 7469 15861 7481 15864
rect 7515 15892 7527 15895
rect 7742 15892 7748 15904
rect 7515 15864 7748 15892
rect 7515 15861 7527 15864
rect 7469 15855 7527 15861
rect 7742 15852 7748 15864
rect 7800 15892 7806 15904
rect 7926 15892 7932 15904
rect 7800 15864 7932 15892
rect 7800 15852 7806 15864
rect 7926 15852 7932 15864
rect 7984 15852 7990 15904
rect 10229 15895 10287 15901
rect 10229 15861 10241 15895
rect 10275 15892 10287 15895
rect 10410 15892 10416 15904
rect 10275 15864 10416 15892
rect 10275 15861 10287 15864
rect 10229 15855 10287 15861
rect 10410 15852 10416 15864
rect 10468 15852 10474 15904
rect 13814 15852 13820 15904
rect 13872 15852 13878 15904
rect 14182 15852 14188 15904
rect 14240 15852 14246 15904
rect 1104 15802 16376 15824
rect 1104 15750 2859 15802
rect 2911 15750 2923 15802
rect 2975 15750 2987 15802
rect 3039 15750 3051 15802
rect 3103 15750 3115 15802
rect 3167 15750 6677 15802
rect 6729 15750 6741 15802
rect 6793 15750 6805 15802
rect 6857 15750 6869 15802
rect 6921 15750 6933 15802
rect 6985 15750 10495 15802
rect 10547 15750 10559 15802
rect 10611 15750 10623 15802
rect 10675 15750 10687 15802
rect 10739 15750 10751 15802
rect 10803 15750 14313 15802
rect 14365 15750 14377 15802
rect 14429 15750 14441 15802
rect 14493 15750 14505 15802
rect 14557 15750 14569 15802
rect 14621 15750 16376 15802
rect 1104 15728 16376 15750
rect 5994 15648 6000 15700
rect 6052 15688 6058 15700
rect 6733 15691 6791 15697
rect 6733 15688 6745 15691
rect 6052 15660 6745 15688
rect 6052 15648 6058 15660
rect 6733 15657 6745 15660
rect 6779 15657 6791 15691
rect 6733 15651 6791 15657
rect 6917 15691 6975 15697
rect 6917 15657 6929 15691
rect 6963 15688 6975 15691
rect 7190 15688 7196 15700
rect 6963 15660 7196 15688
rect 6963 15657 6975 15660
rect 6917 15651 6975 15657
rect 7190 15648 7196 15660
rect 7248 15648 7254 15700
rect 7377 15691 7435 15697
rect 7377 15657 7389 15691
rect 7423 15688 7435 15691
rect 7466 15688 7472 15700
rect 7423 15660 7472 15688
rect 7423 15657 7435 15660
rect 7377 15651 7435 15657
rect 7466 15648 7472 15660
rect 7524 15648 7530 15700
rect 6454 15580 6460 15632
rect 6512 15580 6518 15632
rect 6472 15416 6500 15580
rect 7484 15552 7512 15648
rect 9398 15580 9404 15632
rect 9456 15620 9462 15632
rect 9456 15592 9812 15620
rect 9456 15580 9462 15592
rect 7837 15555 7895 15561
rect 7116 15524 7420 15552
rect 7484 15524 7788 15552
rect 7116 15496 7144 15524
rect 7006 15444 7012 15496
rect 7064 15444 7070 15496
rect 7098 15444 7104 15496
rect 7156 15444 7162 15496
rect 7285 15487 7343 15493
rect 7285 15484 7297 15487
rect 7208 15456 7297 15484
rect 6549 15419 6607 15425
rect 6549 15416 6561 15419
rect 6472 15388 6561 15416
rect 6549 15385 6561 15388
rect 6595 15385 6607 15419
rect 7024 15416 7052 15444
rect 7208 15428 7236 15456
rect 7285 15453 7297 15456
rect 7331 15453 7343 15487
rect 7392 15484 7420 15524
rect 7760 15493 7788 15524
rect 7837 15521 7849 15555
rect 7883 15521 7895 15555
rect 7837 15515 7895 15521
rect 8113 15555 8171 15561
rect 8113 15521 8125 15555
rect 8159 15552 8171 15555
rect 9125 15555 9183 15561
rect 9125 15552 9137 15555
rect 8159 15524 9137 15552
rect 8159 15521 8171 15524
rect 8113 15515 8171 15521
rect 9125 15521 9137 15524
rect 9171 15552 9183 15555
rect 9171 15524 9628 15552
rect 9171 15521 9183 15524
rect 9125 15515 9183 15521
rect 7469 15487 7527 15493
rect 7469 15484 7481 15487
rect 7392 15456 7481 15484
rect 7285 15447 7343 15453
rect 7469 15453 7481 15456
rect 7515 15453 7527 15487
rect 7469 15447 7527 15453
rect 7745 15487 7803 15493
rect 7745 15453 7757 15487
rect 7791 15453 7803 15487
rect 7745 15447 7803 15453
rect 7190 15416 7196 15428
rect 7024 15388 7196 15416
rect 6549 15379 6607 15385
rect 7190 15376 7196 15388
rect 7248 15376 7254 15428
rect 7852 15416 7880 15515
rect 9600 15493 9628 15524
rect 9784 15493 9812 15592
rect 9309 15487 9367 15493
rect 9309 15453 9321 15487
rect 9355 15484 9367 15487
rect 9585 15487 9643 15493
rect 9355 15456 9444 15484
rect 9355 15453 9367 15456
rect 9309 15447 9367 15453
rect 7760 15388 7880 15416
rect 6638 15308 6644 15360
rect 6696 15348 6702 15360
rect 6749 15351 6807 15357
rect 6749 15348 6761 15351
rect 6696 15320 6761 15348
rect 6696 15308 6702 15320
rect 6749 15317 6761 15320
rect 6795 15317 6807 15351
rect 6749 15311 6807 15317
rect 7006 15308 7012 15360
rect 7064 15348 7070 15360
rect 7760 15348 7788 15388
rect 9416 15360 9444 15456
rect 9585 15453 9597 15487
rect 9631 15453 9643 15487
rect 9585 15447 9643 15453
rect 9769 15487 9827 15493
rect 9769 15453 9781 15487
rect 9815 15453 9827 15487
rect 9769 15447 9827 15453
rect 10045 15487 10103 15493
rect 10045 15453 10057 15487
rect 10091 15484 10103 15487
rect 10318 15484 10324 15496
rect 10091 15456 10324 15484
rect 10091 15453 10103 15456
rect 10045 15447 10103 15453
rect 9493 15419 9551 15425
rect 9493 15385 9505 15419
rect 9539 15416 9551 15419
rect 9861 15419 9919 15425
rect 9861 15416 9873 15419
rect 9539 15388 9873 15416
rect 9539 15385 9551 15388
rect 9493 15379 9551 15385
rect 9861 15385 9873 15388
rect 9907 15385 9919 15419
rect 9861 15379 9919 15385
rect 7064 15320 7788 15348
rect 7064 15308 7070 15320
rect 9398 15308 9404 15360
rect 9456 15308 9462 15360
rect 9677 15351 9735 15357
rect 9677 15317 9689 15351
rect 9723 15348 9735 15351
rect 10060 15348 10088 15447
rect 10318 15444 10324 15456
rect 10376 15444 10382 15496
rect 14090 15376 14096 15428
rect 14148 15416 14154 15428
rect 15657 15419 15715 15425
rect 15657 15416 15669 15419
rect 14148 15388 15669 15416
rect 14148 15376 14154 15388
rect 15657 15385 15669 15388
rect 15703 15385 15715 15419
rect 15657 15379 15715 15385
rect 9723 15320 10088 15348
rect 9723 15317 9735 15320
rect 9677 15311 9735 15317
rect 10226 15308 10232 15360
rect 10284 15308 10290 15360
rect 12710 15308 12716 15360
rect 12768 15348 12774 15360
rect 14182 15348 14188 15360
rect 12768 15320 14188 15348
rect 12768 15308 12774 15320
rect 14182 15308 14188 15320
rect 14240 15308 14246 15360
rect 15933 15351 15991 15357
rect 15933 15317 15945 15351
rect 15979 15348 15991 15351
rect 16022 15348 16028 15360
rect 15979 15320 16028 15348
rect 15979 15317 15991 15320
rect 15933 15311 15991 15317
rect 16022 15308 16028 15320
rect 16080 15308 16086 15360
rect 1104 15258 16376 15280
rect 1104 15206 3519 15258
rect 3571 15206 3583 15258
rect 3635 15206 3647 15258
rect 3699 15206 3711 15258
rect 3763 15206 3775 15258
rect 3827 15206 7337 15258
rect 7389 15206 7401 15258
rect 7453 15206 7465 15258
rect 7517 15206 7529 15258
rect 7581 15206 7593 15258
rect 7645 15206 11155 15258
rect 11207 15206 11219 15258
rect 11271 15206 11283 15258
rect 11335 15206 11347 15258
rect 11399 15206 11411 15258
rect 11463 15206 14973 15258
rect 15025 15206 15037 15258
rect 15089 15206 15101 15258
rect 15153 15206 15165 15258
rect 15217 15206 15229 15258
rect 15281 15206 16376 15258
rect 1104 15184 16376 15206
rect 4157 15147 4215 15153
rect 4157 15113 4169 15147
rect 4203 15113 4215 15147
rect 4157 15107 4215 15113
rect 3878 15076 3884 15088
rect 2516 15048 3884 15076
rect 2130 14764 2136 14816
rect 2188 14804 2194 14816
rect 2516 14813 2544 15048
rect 3878 15036 3884 15048
rect 3936 15076 3942 15088
rect 4065 15079 4123 15085
rect 4065 15076 4077 15079
rect 3936 15048 4077 15076
rect 3936 15036 3942 15048
rect 4065 15045 4077 15048
rect 4111 15045 4123 15079
rect 4172 15076 4200 15107
rect 6546 15104 6552 15156
rect 6604 15144 6610 15156
rect 6733 15147 6791 15153
rect 6733 15144 6745 15147
rect 6604 15116 6745 15144
rect 6604 15104 6610 15116
rect 6733 15113 6745 15116
rect 6779 15113 6791 15147
rect 10705 15147 10763 15153
rect 10705 15144 10717 15147
rect 6733 15107 6791 15113
rect 10244 15116 10717 15144
rect 10244 15088 10272 15116
rect 10705 15113 10717 15116
rect 10751 15113 10763 15147
rect 10705 15107 10763 15113
rect 10873 15147 10931 15153
rect 10873 15113 10885 15147
rect 10919 15144 10931 15147
rect 13281 15147 13339 15153
rect 13281 15144 13293 15147
rect 10919 15116 11008 15144
rect 10919 15113 10931 15116
rect 10873 15107 10931 15113
rect 7190 15076 7196 15088
rect 4172 15048 4752 15076
rect 4065 15039 4123 15045
rect 2682 14968 2688 15020
rect 2740 14968 2746 15020
rect 3973 15011 4031 15017
rect 3973 14977 3985 15011
rect 4019 15008 4031 15011
rect 4154 15008 4160 15020
rect 4019 14980 4160 15008
rect 4019 14977 4031 14980
rect 3973 14971 4031 14977
rect 4154 14968 4160 14980
rect 4212 14968 4218 15020
rect 4246 14968 4252 15020
rect 4304 14968 4310 15020
rect 4724 15017 4752 15048
rect 7024 15048 7196 15076
rect 4525 15011 4583 15017
rect 4525 14977 4537 15011
rect 4571 14977 4583 15011
rect 4525 14971 4583 14977
rect 4709 15011 4767 15017
rect 4709 14977 4721 15011
rect 4755 15008 4767 15011
rect 5258 15008 5264 15020
rect 4755 14980 5264 15008
rect 4755 14977 4767 14980
rect 4709 14971 4767 14977
rect 3786 14900 3792 14952
rect 3844 14940 3850 14952
rect 4540 14940 4568 14971
rect 5258 14968 5264 14980
rect 5316 14968 5322 15020
rect 5626 14968 5632 15020
rect 5684 15008 5690 15020
rect 7024 15017 7052 15048
rect 7190 15036 7196 15048
rect 7248 15036 7254 15088
rect 10137 15079 10195 15085
rect 10137 15045 10149 15079
rect 10183 15076 10195 15079
rect 10226 15076 10232 15088
rect 10183 15048 10232 15076
rect 10183 15045 10195 15048
rect 10137 15039 10195 15045
rect 10226 15036 10232 15048
rect 10284 15036 10290 15088
rect 10980 15085 11008 15116
rect 12452 15116 13293 15144
rect 10505 15079 10563 15085
rect 10505 15076 10517 15079
rect 10336 15048 10517 15076
rect 7009 15011 7067 15017
rect 7009 15008 7021 15011
rect 5684 14980 7021 15008
rect 5684 14968 5690 14980
rect 6564 14952 6592 14980
rect 7009 14977 7021 14980
rect 7055 14977 7067 15011
rect 7009 14971 7067 14977
rect 7098 14968 7104 15020
rect 7156 15008 7162 15020
rect 10336 15017 10364 15048
rect 10505 15045 10517 15048
rect 10551 15045 10563 15079
rect 10505 15039 10563 15045
rect 10965 15079 11023 15085
rect 10965 15045 10977 15079
rect 11011 15045 11023 15079
rect 10965 15039 11023 15045
rect 10321 15011 10379 15017
rect 10321 15008 10333 15011
rect 7156 14980 7880 15008
rect 7156 14968 7162 14980
rect 7852 14952 7880 14980
rect 10060 14980 10333 15008
rect 3844 14912 4568 14940
rect 3844 14900 3850 14912
rect 6546 14900 6552 14952
rect 6604 14900 6610 14952
rect 6917 14943 6975 14949
rect 6917 14909 6929 14943
rect 6963 14940 6975 14943
rect 7193 14943 7251 14949
rect 6963 14912 7052 14940
rect 6963 14909 6975 14912
rect 6917 14903 6975 14909
rect 7024 14816 7052 14912
rect 7193 14909 7205 14943
rect 7239 14909 7251 14943
rect 7193 14903 7251 14909
rect 7208 14816 7236 14903
rect 7834 14900 7840 14952
rect 7892 14900 7898 14952
rect 10060 14816 10088 14980
rect 10321 14977 10333 14980
rect 10367 14977 10379 15011
rect 10321 14971 10379 14977
rect 10413 15011 10471 15017
rect 10413 14977 10425 15011
rect 10459 15008 10471 15011
rect 10594 15008 10600 15020
rect 10459 14980 10600 15008
rect 10459 14977 10471 14980
rect 10413 14971 10471 14977
rect 10594 14968 10600 14980
rect 10652 14968 10658 15020
rect 12452 15017 12480 15116
rect 13281 15113 13293 15116
rect 13327 15113 13339 15147
rect 13281 15107 13339 15113
rect 12529 15079 12587 15085
rect 12529 15045 12541 15079
rect 12575 15076 12587 15079
rect 12710 15076 12716 15088
rect 12575 15048 12716 15076
rect 12575 15045 12587 15048
rect 12529 15039 12587 15045
rect 12710 15036 12716 15048
rect 12768 15036 12774 15088
rect 13081 15079 13139 15085
rect 13081 15076 13093 15079
rect 12820 15048 13093 15076
rect 12820 15017 12848 15048
rect 13081 15045 13093 15048
rect 13127 15045 13139 15079
rect 14277 15079 14335 15085
rect 14277 15076 14289 15079
rect 13081 15039 13139 15045
rect 14016 15048 14289 15076
rect 11149 15011 11207 15017
rect 11149 14977 11161 15011
rect 11195 14977 11207 15011
rect 11149 14971 11207 14977
rect 12437 15011 12495 15017
rect 12437 14977 12449 15011
rect 12483 14977 12495 15011
rect 12437 14971 12495 14977
rect 12805 15011 12863 15017
rect 12805 14977 12817 15011
rect 12851 14977 12863 15011
rect 12805 14971 12863 14977
rect 13725 15011 13783 15017
rect 13725 14977 13737 15011
rect 13771 15008 13783 15011
rect 13906 15008 13912 15020
rect 13771 14980 13912 15008
rect 13771 14977 13783 14980
rect 13725 14971 13783 14977
rect 11164 14940 11192 14971
rect 10520 14912 11192 14940
rect 11333 14943 11391 14949
rect 2501 14807 2559 14813
rect 2501 14804 2513 14807
rect 2188 14776 2513 14804
rect 2188 14764 2194 14776
rect 2501 14773 2513 14776
rect 2547 14773 2559 14807
rect 2501 14767 2559 14773
rect 4617 14807 4675 14813
rect 4617 14773 4629 14807
rect 4663 14804 4675 14807
rect 5166 14804 5172 14816
rect 4663 14776 5172 14804
rect 4663 14773 4675 14776
rect 4617 14767 4675 14773
rect 5166 14764 5172 14776
rect 5224 14764 5230 14816
rect 7006 14764 7012 14816
rect 7064 14764 7070 14816
rect 7190 14764 7196 14816
rect 7248 14764 7254 14816
rect 10042 14764 10048 14816
rect 10100 14764 10106 14816
rect 10134 14764 10140 14816
rect 10192 14804 10198 14816
rect 10520 14804 10548 14912
rect 11333 14909 11345 14943
rect 11379 14940 11391 14943
rect 12452 14940 12480 14971
rect 11379 14912 12480 14940
rect 11379 14909 11391 14912
rect 11333 14903 11391 14909
rect 12820 14816 12848 14971
rect 13906 14968 13912 14980
rect 13964 14968 13970 15020
rect 12989 14943 13047 14949
rect 12989 14909 13001 14943
rect 13035 14909 13047 14943
rect 12989 14903 13047 14909
rect 13004 14816 13032 14903
rect 13814 14900 13820 14952
rect 13872 14940 13878 14952
rect 14016 14940 14044 15048
rect 14277 15045 14289 15048
rect 14323 15045 14335 15079
rect 14277 15039 14335 15045
rect 14182 14968 14188 15020
rect 14240 14968 14246 15020
rect 14369 15011 14427 15017
rect 14369 15008 14381 15011
rect 14292 14980 14381 15008
rect 13872 14912 14044 14940
rect 13872 14900 13878 14912
rect 14090 14900 14096 14952
rect 14148 14900 14154 14952
rect 13449 14875 13507 14881
rect 13449 14841 13461 14875
rect 13495 14872 13507 14875
rect 14292 14872 14320 14980
rect 14369 14977 14381 14980
rect 14415 14977 14427 15011
rect 14369 14971 14427 14977
rect 13495 14844 14320 14872
rect 13495 14841 13507 14844
rect 13449 14835 13507 14841
rect 10192 14776 10548 14804
rect 10192 14764 10198 14776
rect 10594 14764 10600 14816
rect 10652 14804 10658 14816
rect 10689 14807 10747 14813
rect 10689 14804 10701 14807
rect 10652 14776 10701 14804
rect 10652 14764 10658 14776
rect 10689 14773 10701 14776
rect 10735 14804 10747 14807
rect 10962 14804 10968 14816
rect 10735 14776 10968 14804
rect 10735 14773 10747 14776
rect 10689 14767 10747 14773
rect 10962 14764 10968 14776
rect 11020 14764 11026 14816
rect 12802 14764 12808 14816
rect 12860 14764 12866 14816
rect 12986 14764 12992 14816
rect 13044 14804 13050 14816
rect 13265 14807 13323 14813
rect 13265 14804 13277 14807
rect 13044 14776 13277 14804
rect 13044 14764 13050 14776
rect 13265 14773 13277 14776
rect 13311 14773 13323 14807
rect 13265 14767 13323 14773
rect 1104 14714 16376 14736
rect 1104 14662 2859 14714
rect 2911 14662 2923 14714
rect 2975 14662 2987 14714
rect 3039 14662 3051 14714
rect 3103 14662 3115 14714
rect 3167 14662 6677 14714
rect 6729 14662 6741 14714
rect 6793 14662 6805 14714
rect 6857 14662 6869 14714
rect 6921 14662 6933 14714
rect 6985 14662 10495 14714
rect 10547 14662 10559 14714
rect 10611 14662 10623 14714
rect 10675 14662 10687 14714
rect 10739 14662 10751 14714
rect 10803 14662 14313 14714
rect 14365 14662 14377 14714
rect 14429 14662 14441 14714
rect 14493 14662 14505 14714
rect 14557 14662 14569 14714
rect 14621 14662 16376 14714
rect 1104 14640 16376 14662
rect 4062 14600 4068 14612
rect 2608 14572 4068 14600
rect 2501 14399 2559 14405
rect 2501 14365 2513 14399
rect 2547 14396 2559 14399
rect 2608 14396 2636 14572
rect 4062 14560 4068 14572
rect 4120 14560 4126 14612
rect 4617 14603 4675 14609
rect 4617 14600 4629 14603
rect 4172 14572 4629 14600
rect 3326 14492 3332 14544
rect 3384 14492 3390 14544
rect 4172 14532 4200 14572
rect 4617 14569 4629 14572
rect 4663 14569 4675 14603
rect 4617 14563 4675 14569
rect 3620 14504 4200 14532
rect 4433 14535 4491 14541
rect 3510 14464 3516 14476
rect 3344 14436 3516 14464
rect 2547 14368 2636 14396
rect 2685 14399 2743 14405
rect 2547 14365 2559 14368
rect 2501 14359 2559 14365
rect 2685 14365 2697 14399
rect 2731 14365 2743 14399
rect 2685 14359 2743 14365
rect 2869 14399 2927 14405
rect 2869 14365 2881 14399
rect 2915 14365 2927 14399
rect 2869 14359 2927 14365
rect 934 14288 940 14340
rect 992 14328 998 14340
rect 1489 14331 1547 14337
rect 1489 14328 1501 14331
rect 992 14300 1501 14328
rect 992 14288 998 14300
rect 1489 14297 1501 14300
rect 1535 14297 1547 14331
rect 1489 14291 1547 14297
rect 2590 14288 2596 14340
rect 2648 14328 2654 14340
rect 2700 14328 2728 14359
rect 2648 14300 2728 14328
rect 2648 14288 2654 14300
rect 2774 14288 2780 14340
rect 2832 14288 2838 14340
rect 1394 14220 1400 14272
rect 1452 14260 1458 14272
rect 1581 14263 1639 14269
rect 1581 14260 1593 14263
rect 1452 14232 1593 14260
rect 1452 14220 1458 14232
rect 1581 14229 1593 14232
rect 1627 14260 1639 14263
rect 2222 14260 2228 14272
rect 1627 14232 2228 14260
rect 1627 14229 1639 14232
rect 1581 14223 1639 14229
rect 2222 14220 2228 14232
rect 2280 14260 2286 14272
rect 2682 14260 2688 14272
rect 2280 14232 2688 14260
rect 2280 14220 2286 14232
rect 2682 14220 2688 14232
rect 2740 14260 2746 14272
rect 2884 14260 2912 14359
rect 3234 14356 3240 14408
rect 3292 14396 3298 14408
rect 3344 14405 3372 14436
rect 3510 14424 3516 14436
rect 3568 14424 3574 14476
rect 3620 14405 3648 14504
rect 4433 14501 4445 14535
rect 4479 14501 4491 14535
rect 4433 14495 4491 14501
rect 3786 14424 3792 14476
rect 3844 14424 3850 14476
rect 3878 14424 3884 14476
rect 3936 14464 3942 14476
rect 4065 14467 4123 14473
rect 4065 14464 4077 14467
rect 3936 14436 4077 14464
rect 3936 14424 3942 14436
rect 4065 14433 4077 14436
rect 4111 14433 4123 14467
rect 4065 14427 4123 14433
rect 4246 14424 4252 14476
rect 4304 14464 4310 14476
rect 4448 14464 4476 14495
rect 4304 14436 4476 14464
rect 4632 14464 4660 14563
rect 5258 14560 5264 14612
rect 5316 14600 5322 14612
rect 5629 14603 5687 14609
rect 5629 14600 5641 14603
rect 5316 14572 5641 14600
rect 5316 14560 5322 14572
rect 5629 14569 5641 14572
rect 5675 14569 5687 14603
rect 5629 14563 5687 14569
rect 9398 14560 9404 14612
rect 9456 14560 9462 14612
rect 10042 14560 10048 14612
rect 10100 14560 10106 14612
rect 10962 14560 10968 14612
rect 11020 14560 11026 14612
rect 12437 14603 12495 14609
rect 12437 14569 12449 14603
rect 12483 14569 12495 14603
rect 12437 14563 12495 14569
rect 5813 14535 5871 14541
rect 5813 14501 5825 14535
rect 5859 14532 5871 14535
rect 5859 14504 10088 14532
rect 5859 14501 5871 14504
rect 5813 14495 5871 14501
rect 5997 14467 6055 14473
rect 4632 14436 5488 14464
rect 4304 14424 4310 14436
rect 3329 14399 3387 14405
rect 3329 14396 3341 14399
rect 3292 14368 3341 14396
rect 3292 14356 3298 14368
rect 3329 14365 3341 14368
rect 3375 14365 3387 14399
rect 3605 14399 3663 14405
rect 3605 14396 3617 14399
rect 3329 14359 3387 14365
rect 3436 14368 3617 14396
rect 3436 14340 3464 14368
rect 3605 14365 3617 14368
rect 3651 14365 3663 14399
rect 3605 14359 3663 14365
rect 3970 14356 3976 14408
rect 4028 14356 4034 14408
rect 4154 14356 4160 14408
rect 4212 14396 4218 14408
rect 4522 14396 4528 14408
rect 4212 14368 4528 14396
rect 4212 14356 4218 14368
rect 4522 14356 4528 14368
rect 4580 14356 4586 14408
rect 4893 14399 4951 14405
rect 4893 14365 4905 14399
rect 4939 14396 4951 14399
rect 4939 14368 5120 14396
rect 4939 14365 4951 14368
rect 4893 14359 4951 14365
rect 3418 14288 3424 14340
rect 3476 14288 3482 14340
rect 3513 14331 3571 14337
rect 3513 14297 3525 14331
rect 3559 14328 3571 14331
rect 4801 14331 4859 14337
rect 4801 14328 4813 14331
rect 3559 14300 4813 14328
rect 3559 14297 3571 14300
rect 3513 14291 3571 14297
rect 4801 14297 4813 14300
rect 4847 14297 4859 14331
rect 4801 14291 4859 14297
rect 2740 14232 2912 14260
rect 3053 14263 3111 14269
rect 2740 14220 2746 14232
rect 3053 14229 3065 14263
rect 3099 14260 3111 14263
rect 3528 14260 3556 14291
rect 5092 14272 5120 14368
rect 5166 14356 5172 14408
rect 5224 14356 5230 14408
rect 5460 14337 5488 14436
rect 5997 14433 6009 14467
rect 6043 14464 6055 14467
rect 6043 14436 8800 14464
rect 6043 14433 6055 14436
rect 5997 14427 6055 14433
rect 5902 14356 5908 14408
rect 5960 14356 5966 14408
rect 6089 14399 6147 14405
rect 6089 14365 6101 14399
rect 6135 14365 6147 14399
rect 6089 14359 6147 14365
rect 5445 14331 5503 14337
rect 5445 14297 5457 14331
rect 5491 14297 5503 14331
rect 6104 14328 6132 14359
rect 7190 14328 7196 14340
rect 5445 14291 5503 14297
rect 5736 14300 6132 14328
rect 6748 14300 7196 14328
rect 3099 14232 3556 14260
rect 3099 14229 3111 14232
rect 3053 14223 3111 14229
rect 3602 14220 3608 14272
rect 3660 14260 3666 14272
rect 4591 14263 4649 14269
rect 4591 14260 4603 14263
rect 3660 14232 4603 14260
rect 3660 14220 3666 14232
rect 4591 14229 4603 14232
rect 4637 14229 4649 14263
rect 4591 14223 4649 14229
rect 4982 14220 4988 14272
rect 5040 14220 5046 14272
rect 5074 14220 5080 14272
rect 5132 14220 5138 14272
rect 5353 14263 5411 14269
rect 5353 14229 5365 14263
rect 5399 14260 5411 14263
rect 5645 14263 5703 14269
rect 5645 14260 5657 14263
rect 5399 14232 5657 14260
rect 5399 14229 5411 14232
rect 5353 14223 5411 14229
rect 5645 14229 5657 14232
rect 5691 14260 5703 14263
rect 5736 14260 5764 14300
rect 6748 14272 6776 14300
rect 7190 14288 7196 14300
rect 7248 14288 7254 14340
rect 7377 14331 7435 14337
rect 7377 14297 7389 14331
rect 7423 14328 7435 14331
rect 8018 14328 8024 14340
rect 7423 14300 8024 14328
rect 7423 14297 7435 14300
rect 7377 14291 7435 14297
rect 8018 14288 8024 14300
rect 8076 14288 8082 14340
rect 8772 14328 8800 14436
rect 8846 14424 8852 14476
rect 8904 14464 8910 14476
rect 9033 14467 9091 14473
rect 9033 14464 9045 14467
rect 8904 14436 9045 14464
rect 8904 14424 8910 14436
rect 9033 14433 9045 14436
rect 9079 14433 9091 14467
rect 9033 14427 9091 14433
rect 9125 14399 9183 14405
rect 9125 14365 9137 14399
rect 9171 14396 9183 14399
rect 9214 14396 9220 14408
rect 9171 14368 9220 14396
rect 9171 14365 9183 14368
rect 9125 14359 9183 14365
rect 9214 14356 9220 14368
rect 9272 14356 9278 14408
rect 10060 14396 10088 14504
rect 10980 14464 11008 14560
rect 12452 14532 12480 14563
rect 12802 14560 12808 14612
rect 12860 14560 12866 14612
rect 12406 14504 12480 14532
rect 11057 14467 11115 14473
rect 11057 14464 11069 14467
rect 10980 14436 11069 14464
rect 11057 14433 11069 14436
rect 11103 14433 11115 14467
rect 11793 14467 11851 14473
rect 11793 14464 11805 14467
rect 11057 14427 11115 14433
rect 11164 14436 11805 14464
rect 11164 14396 11192 14436
rect 11793 14433 11805 14436
rect 11839 14464 11851 14467
rect 12406 14464 12434 14504
rect 11839 14436 12434 14464
rect 11839 14433 11851 14436
rect 11793 14427 11851 14433
rect 9600 14368 9996 14396
rect 10060 14368 11192 14396
rect 11241 14399 11299 14405
rect 9600 14328 9628 14368
rect 8772 14300 9628 14328
rect 9674 14288 9680 14340
rect 9732 14288 9738 14340
rect 9861 14331 9919 14337
rect 9861 14297 9873 14331
rect 9907 14297 9919 14331
rect 9861 14291 9919 14297
rect 5691 14232 5764 14260
rect 5691 14229 5703 14232
rect 5645 14223 5703 14229
rect 6730 14220 6736 14272
rect 6788 14220 6794 14272
rect 7561 14263 7619 14269
rect 7561 14229 7573 14263
rect 7607 14260 7619 14263
rect 9766 14260 9772 14272
rect 7607 14232 9772 14260
rect 7607 14229 7619 14232
rect 7561 14223 7619 14229
rect 9766 14220 9772 14232
rect 9824 14260 9830 14272
rect 9876 14260 9904 14291
rect 9824 14232 9904 14260
rect 9968 14260 9996 14368
rect 11241 14365 11253 14399
rect 11287 14365 11299 14399
rect 11241 14359 11299 14365
rect 11425 14399 11483 14405
rect 11425 14365 11437 14399
rect 11471 14396 11483 14399
rect 11885 14399 11943 14405
rect 11885 14396 11897 14399
rect 11471 14368 11897 14396
rect 11471 14365 11483 14368
rect 11425 14359 11483 14365
rect 11885 14365 11897 14368
rect 11931 14396 11943 14399
rect 12345 14399 12403 14405
rect 12345 14396 12357 14399
rect 11931 14368 12357 14396
rect 11931 14365 11943 14368
rect 11885 14359 11943 14365
rect 12345 14365 12357 14368
rect 12391 14365 12403 14399
rect 12345 14359 12403 14365
rect 10594 14288 10600 14340
rect 10652 14288 10658 14340
rect 10778 14288 10784 14340
rect 10836 14288 10842 14340
rect 10870 14288 10876 14340
rect 10928 14328 10934 14340
rect 11256 14328 11284 14359
rect 10928 14300 11284 14328
rect 10928 14288 10934 14300
rect 11054 14260 11060 14272
rect 9968 14232 11060 14260
rect 9824 14220 9830 14232
rect 11054 14220 11060 14232
rect 11112 14220 11118 14272
rect 12253 14263 12311 14269
rect 12253 14229 12265 14263
rect 12299 14260 12311 14263
rect 12710 14260 12716 14272
rect 12299 14232 12716 14260
rect 12299 14229 12311 14232
rect 12253 14223 12311 14229
rect 12710 14220 12716 14232
rect 12768 14220 12774 14272
rect 1104 14170 16376 14192
rect 1104 14118 3519 14170
rect 3571 14118 3583 14170
rect 3635 14118 3647 14170
rect 3699 14118 3711 14170
rect 3763 14118 3775 14170
rect 3827 14118 7337 14170
rect 7389 14118 7401 14170
rect 7453 14118 7465 14170
rect 7517 14118 7529 14170
rect 7581 14118 7593 14170
rect 7645 14118 11155 14170
rect 11207 14118 11219 14170
rect 11271 14118 11283 14170
rect 11335 14118 11347 14170
rect 11399 14118 11411 14170
rect 11463 14118 14973 14170
rect 15025 14118 15037 14170
rect 15089 14118 15101 14170
rect 15153 14118 15165 14170
rect 15217 14118 15229 14170
rect 15281 14118 16376 14170
rect 1104 14096 16376 14118
rect 1946 14056 1952 14068
rect 1596 14028 1952 14056
rect 1394 13948 1400 14000
rect 1452 13948 1458 14000
rect 1596 13997 1624 14028
rect 1946 14016 1952 14028
rect 2004 14016 2010 14068
rect 2222 14016 2228 14068
rect 2280 14056 2286 14068
rect 2685 14059 2743 14065
rect 2280 14028 2636 14056
rect 2280 14016 2286 14028
rect 1581 13991 1639 13997
rect 1581 13957 1593 13991
rect 1627 13957 1639 13991
rect 1581 13951 1639 13957
rect 1673 13991 1731 13997
rect 1673 13957 1685 13991
rect 1719 13988 1731 13991
rect 2317 13991 2375 13997
rect 2317 13988 2329 13991
rect 1719 13960 2329 13988
rect 1719 13957 1731 13960
rect 1673 13951 1731 13957
rect 2317 13957 2329 13960
rect 2363 13988 2375 13991
rect 2498 13988 2504 14000
rect 2363 13960 2504 13988
rect 2363 13957 2375 13960
rect 2317 13951 2375 13957
rect 2498 13948 2504 13960
rect 2556 13948 2562 14000
rect 2608 13988 2636 14028
rect 2685 14025 2697 14059
rect 2731 14056 2743 14059
rect 3234 14056 3240 14068
rect 2731 14028 3240 14056
rect 2731 14025 2743 14028
rect 2685 14019 2743 14025
rect 3234 14016 3240 14028
rect 3292 14016 3298 14068
rect 3418 14016 3424 14068
rect 3476 14056 3482 14068
rect 3605 14059 3663 14065
rect 3605 14056 3617 14059
rect 3476 14028 3617 14056
rect 3476 14016 3482 14028
rect 3605 14025 3617 14028
rect 3651 14025 3663 14059
rect 3605 14019 3663 14025
rect 3970 14016 3976 14068
rect 4028 14016 4034 14068
rect 5166 14016 5172 14068
rect 5224 14016 5230 14068
rect 5261 14059 5319 14065
rect 5261 14025 5273 14059
rect 5307 14056 5319 14059
rect 5902 14056 5908 14068
rect 5307 14028 5908 14056
rect 5307 14025 5319 14028
rect 5261 14019 5319 14025
rect 5902 14016 5908 14028
rect 5960 14016 5966 14068
rect 6730 14016 6736 14068
rect 6788 14016 6794 14068
rect 7009 14059 7067 14065
rect 7009 14025 7021 14059
rect 7055 14056 7067 14059
rect 7282 14056 7288 14068
rect 7055 14028 7288 14056
rect 7055 14025 7067 14028
rect 7009 14019 7067 14025
rect 7282 14016 7288 14028
rect 7340 14056 7346 14068
rect 7742 14056 7748 14068
rect 7340 14028 7748 14056
rect 7340 14016 7346 14028
rect 7742 14016 7748 14028
rect 7800 14016 7806 14068
rect 8938 14016 8944 14068
rect 8996 14016 9002 14068
rect 9401 14059 9459 14065
rect 9401 14025 9413 14059
rect 9447 14056 9459 14059
rect 9674 14056 9680 14068
rect 9447 14028 9680 14056
rect 9447 14025 9459 14028
rect 9401 14019 9459 14025
rect 3988 13988 4016 14016
rect 2608 13960 3004 13988
rect 1412 13920 1440 13948
rect 1484 13929 1542 13935
rect 1484 13920 1496 13929
rect 1412 13895 1496 13920
rect 1530 13895 1542 13929
rect 1412 13892 1542 13895
rect 1484 13889 1542 13892
rect 1857 13923 1915 13929
rect 1857 13889 1869 13923
rect 1903 13920 1915 13923
rect 1903 13892 2176 13920
rect 1903 13889 1915 13892
rect 1857 13883 1915 13889
rect 1872 13784 1900 13883
rect 1946 13812 1952 13864
rect 2004 13812 2010 13864
rect 2148 13852 2176 13892
rect 2222 13880 2228 13932
rect 2280 13880 2286 13932
rect 2976 13929 3004 13960
rect 3252 13960 4016 13988
rect 4985 13991 5043 13997
rect 3252 13929 3280 13960
rect 4985 13957 4997 13991
rect 5031 13988 5043 13991
rect 5184 13988 5212 14016
rect 5031 13960 5212 13988
rect 5031 13957 5043 13960
rect 4985 13951 5043 13957
rect 7190 13948 7196 14000
rect 7248 13988 7254 14000
rect 7423 13991 7481 13997
rect 7423 13988 7435 13991
rect 7248 13960 7435 13988
rect 7248 13948 7254 13960
rect 7423 13957 7435 13960
rect 7469 13957 7481 13991
rect 7423 13951 7481 13957
rect 7760 13951 7788 14016
rect 9214 13988 9220 14000
rect 8680 13960 9220 13988
rect 7750 13945 7808 13951
rect 2409 13923 2467 13929
rect 2409 13889 2421 13923
rect 2455 13889 2467 13923
rect 2409 13883 2467 13889
rect 2961 13923 3019 13929
rect 2961 13889 2973 13923
rect 3007 13889 3019 13923
rect 2961 13883 3019 13889
rect 3237 13923 3295 13929
rect 3237 13889 3249 13923
rect 3283 13889 3295 13923
rect 3237 13883 3295 13889
rect 2424 13852 2452 13883
rect 2148 13824 2452 13852
rect 2682 13812 2688 13864
rect 2740 13852 2746 13864
rect 3252 13852 3280 13883
rect 3418 13880 3424 13932
rect 3476 13920 3482 13932
rect 4157 13923 4215 13929
rect 4157 13920 4169 13923
rect 3476 13892 4169 13920
rect 3476 13880 3482 13892
rect 4157 13889 4169 13892
rect 4203 13889 4215 13923
rect 4157 13883 4215 13889
rect 4246 13880 4252 13932
rect 4304 13920 4310 13932
rect 4341 13923 4399 13929
rect 4341 13920 4353 13923
rect 4304 13892 4353 13920
rect 4304 13880 4310 13892
rect 4341 13889 4353 13892
rect 4387 13889 4399 13923
rect 4341 13883 4399 13889
rect 5074 13880 5080 13932
rect 5132 13920 5138 13932
rect 5169 13923 5227 13929
rect 5169 13920 5181 13923
rect 5132 13892 5181 13920
rect 5132 13880 5138 13892
rect 5169 13889 5181 13892
rect 5215 13889 5227 13923
rect 5169 13883 5227 13889
rect 5261 13923 5319 13929
rect 5261 13889 5273 13923
rect 5307 13920 5319 13923
rect 6917 13923 6975 13929
rect 5307 13892 5396 13920
rect 5307 13889 5319 13892
rect 5261 13883 5319 13889
rect 5368 13864 5396 13892
rect 6917 13889 6929 13923
rect 6963 13889 6975 13923
rect 6917 13883 6975 13889
rect 2740 13824 3280 13852
rect 3329 13855 3387 13861
rect 2740 13812 2746 13824
rect 3329 13821 3341 13855
rect 3375 13852 3387 13855
rect 3375 13824 4936 13852
rect 3375 13821 3387 13824
rect 3329 13815 3387 13821
rect 2041 13787 2099 13793
rect 1872 13756 1992 13784
rect 1964 13728 1992 13756
rect 2041 13753 2053 13787
rect 2087 13784 2099 13787
rect 2774 13784 2780 13796
rect 2087 13756 2780 13784
rect 2087 13753 2099 13756
rect 2041 13747 2099 13753
rect 2774 13744 2780 13756
rect 2832 13744 2838 13796
rect 1854 13676 1860 13728
rect 1912 13676 1918 13728
rect 1946 13676 1952 13728
rect 2004 13676 2010 13728
rect 3053 13719 3111 13725
rect 3053 13685 3065 13719
rect 3099 13716 3111 13719
rect 3237 13719 3295 13725
rect 3237 13716 3249 13719
rect 3099 13688 3249 13716
rect 3099 13685 3111 13688
rect 3053 13679 3111 13685
rect 3237 13685 3249 13688
rect 3283 13685 3295 13719
rect 3237 13679 3295 13685
rect 4154 13676 4160 13728
rect 4212 13676 4218 13728
rect 4908 13716 4936 13824
rect 4982 13812 4988 13864
rect 5040 13852 5046 13864
rect 5350 13852 5356 13864
rect 5040 13824 5356 13852
rect 5040 13812 5046 13824
rect 5350 13812 5356 13824
rect 5408 13812 5414 13864
rect 6932 13852 6960 13883
rect 7098 13880 7104 13932
rect 7156 13880 7162 13932
rect 7558 13920 7564 13932
rect 7192 13892 7564 13920
rect 7192 13852 7220 13892
rect 7558 13880 7564 13892
rect 7616 13880 7622 13932
rect 7650 13880 7656 13932
rect 7708 13880 7714 13932
rect 7750 13911 7762 13945
rect 7796 13911 7808 13945
rect 7750 13905 7808 13911
rect 6932 13824 7220 13852
rect 7469 13855 7527 13861
rect 5258 13744 5264 13796
rect 5316 13784 5322 13796
rect 6546 13784 6552 13796
rect 5316 13756 6552 13784
rect 5316 13744 5322 13756
rect 6546 13744 6552 13756
rect 6604 13784 6610 13796
rect 6932 13784 6960 13824
rect 7469 13821 7481 13855
rect 7515 13852 7527 13855
rect 8018 13852 8024 13864
rect 7515 13824 7604 13852
rect 7515 13821 7527 13824
rect 7469 13815 7527 13821
rect 6604 13756 6960 13784
rect 6604 13744 6610 13756
rect 7190 13744 7196 13796
rect 7248 13784 7254 13796
rect 7285 13787 7343 13793
rect 7285 13784 7297 13787
rect 7248 13756 7297 13784
rect 7248 13744 7254 13756
rect 7285 13753 7297 13756
rect 7331 13753 7343 13787
rect 7576 13784 7604 13824
rect 7852 13824 8024 13852
rect 7852 13784 7880 13824
rect 8018 13812 8024 13824
rect 8076 13812 8082 13864
rect 8297 13855 8355 13861
rect 8297 13821 8309 13855
rect 8343 13852 8355 13855
rect 8386 13852 8392 13864
rect 8343 13824 8392 13852
rect 8343 13821 8355 13824
rect 8297 13815 8355 13821
rect 8386 13812 8392 13824
rect 8444 13812 8450 13864
rect 8570 13812 8576 13864
rect 8628 13852 8634 13864
rect 8680 13861 8708 13960
rect 9214 13948 9220 13960
rect 9272 13948 9278 14000
rect 9033 13923 9091 13929
rect 9033 13889 9045 13923
rect 9079 13920 9091 13923
rect 9122 13920 9128 13932
rect 9079 13892 9128 13920
rect 9079 13889 9091 13892
rect 9033 13883 9091 13889
rect 9122 13880 9128 13892
rect 9180 13880 9186 13932
rect 8665 13855 8723 13861
rect 8665 13852 8677 13855
rect 8628 13824 8677 13852
rect 8628 13812 8634 13824
rect 8665 13821 8677 13824
rect 8711 13821 8723 13855
rect 8665 13815 8723 13821
rect 8757 13855 8815 13861
rect 8757 13821 8769 13855
rect 8803 13852 8815 13855
rect 8846 13852 8852 13864
rect 8803 13824 8852 13852
rect 8803 13821 8815 13824
rect 8757 13815 8815 13821
rect 8846 13812 8852 13824
rect 8904 13812 8910 13864
rect 9600 13861 9628 14028
rect 9674 14016 9680 14028
rect 9732 14016 9738 14068
rect 9766 14016 9772 14068
rect 9824 14016 9830 14068
rect 10870 14016 10876 14068
rect 10928 14016 10934 14068
rect 9677 13923 9735 13929
rect 9677 13889 9689 13923
rect 9723 13920 9735 13923
rect 9784 13920 9812 14016
rect 10594 13920 10600 13932
rect 9723 13892 9812 13920
rect 10060 13892 10600 13920
rect 9723 13889 9735 13892
rect 9677 13883 9735 13889
rect 9585 13855 9643 13861
rect 9585 13821 9597 13855
rect 9631 13821 9643 13855
rect 9585 13815 9643 13821
rect 10060 13793 10088 13892
rect 10594 13880 10600 13892
rect 10652 13920 10658 13932
rect 10689 13923 10747 13929
rect 10689 13920 10701 13923
rect 10652 13892 10701 13920
rect 10652 13880 10658 13892
rect 10689 13889 10701 13892
rect 10735 13889 10747 13923
rect 10689 13883 10747 13889
rect 10870 13880 10876 13932
rect 10928 13880 10934 13932
rect 7576 13756 7880 13784
rect 10045 13787 10103 13793
rect 7285 13747 7343 13753
rect 10045 13753 10057 13787
rect 10091 13753 10103 13787
rect 10045 13747 10103 13753
rect 5994 13716 6000 13728
rect 4908 13688 6000 13716
rect 5994 13676 6000 13688
rect 6052 13676 6058 13728
rect 1104 13626 16376 13648
rect 1104 13574 2859 13626
rect 2911 13574 2923 13626
rect 2975 13574 2987 13626
rect 3039 13574 3051 13626
rect 3103 13574 3115 13626
rect 3167 13574 6677 13626
rect 6729 13574 6741 13626
rect 6793 13574 6805 13626
rect 6857 13574 6869 13626
rect 6921 13574 6933 13626
rect 6985 13574 10495 13626
rect 10547 13574 10559 13626
rect 10611 13574 10623 13626
rect 10675 13574 10687 13626
rect 10739 13574 10751 13626
rect 10803 13574 14313 13626
rect 14365 13574 14377 13626
rect 14429 13574 14441 13626
rect 14493 13574 14505 13626
rect 14557 13574 14569 13626
rect 14621 13574 16376 13626
rect 1104 13552 16376 13574
rect 2590 13472 2596 13524
rect 2648 13472 2654 13524
rect 2774 13472 2780 13524
rect 2832 13512 2838 13524
rect 3053 13515 3111 13521
rect 3053 13512 3065 13515
rect 2832 13484 3065 13512
rect 2832 13472 2838 13484
rect 3053 13481 3065 13484
rect 3099 13481 3111 13515
rect 3513 13515 3571 13521
rect 3513 13512 3525 13515
rect 3053 13475 3111 13481
rect 3160 13484 3525 13512
rect 2608 13444 2636 13472
rect 3160 13444 3188 13484
rect 3513 13481 3525 13484
rect 3559 13512 3571 13515
rect 5258 13512 5264 13524
rect 3559 13484 5264 13512
rect 3559 13481 3571 13484
rect 3513 13475 3571 13481
rect 5258 13472 5264 13484
rect 5316 13472 5322 13524
rect 5350 13472 5356 13524
rect 5408 13512 5414 13524
rect 5905 13515 5963 13521
rect 5905 13512 5917 13515
rect 5408 13484 5917 13512
rect 5408 13472 5414 13484
rect 5905 13481 5917 13484
rect 5951 13481 5963 13515
rect 5905 13475 5963 13481
rect 7006 13472 7012 13524
rect 7064 13472 7070 13524
rect 7193 13515 7251 13521
rect 7193 13481 7205 13515
rect 7239 13512 7251 13515
rect 7282 13512 7288 13524
rect 7239 13484 7288 13512
rect 7239 13481 7251 13484
rect 7193 13475 7251 13481
rect 7282 13472 7288 13484
rect 7340 13472 7346 13524
rect 7558 13472 7564 13524
rect 7616 13472 7622 13524
rect 8386 13472 8392 13524
rect 8444 13472 8450 13524
rect 8570 13472 8576 13524
rect 8628 13472 8634 13524
rect 9122 13472 9128 13524
rect 9180 13512 9186 13524
rect 9217 13515 9275 13521
rect 9217 13512 9229 13515
rect 9180 13484 9229 13512
rect 9180 13472 9186 13484
rect 9217 13481 9229 13484
rect 9263 13481 9275 13515
rect 9217 13475 9275 13481
rect 12342 13472 12348 13524
rect 12400 13512 12406 13524
rect 12805 13515 12863 13521
rect 12805 13512 12817 13515
rect 12400 13484 12817 13512
rect 12400 13472 12406 13484
rect 12805 13481 12817 13484
rect 12851 13481 12863 13515
rect 12805 13475 12863 13481
rect 12986 13472 12992 13524
rect 13044 13472 13050 13524
rect 13906 13472 13912 13524
rect 13964 13512 13970 13524
rect 14093 13515 14151 13521
rect 14093 13512 14105 13515
rect 13964 13484 14105 13512
rect 13964 13472 13970 13484
rect 14093 13481 14105 13484
rect 14139 13481 14151 13515
rect 14093 13475 14151 13481
rect 2608 13416 3188 13444
rect 3252 13416 6500 13444
rect 1854 13336 1860 13388
rect 1912 13376 1918 13388
rect 1949 13379 2007 13385
rect 1949 13376 1961 13379
rect 1912 13348 1961 13376
rect 1912 13336 1918 13348
rect 1949 13345 1961 13348
rect 1995 13345 2007 13379
rect 1949 13339 2007 13345
rect 2130 13336 2136 13388
rect 2188 13336 2194 13388
rect 3252 13320 3280 13416
rect 5276 13348 5948 13376
rect 934 13268 940 13320
rect 992 13308 998 13320
rect 1397 13311 1455 13317
rect 1397 13308 1409 13311
rect 992 13280 1409 13308
rect 992 13268 998 13280
rect 1397 13277 1409 13280
rect 1443 13277 1455 13311
rect 1397 13271 1455 13277
rect 2041 13311 2099 13317
rect 2041 13277 2053 13311
rect 2087 13277 2099 13311
rect 2041 13271 2099 13277
rect 1946 13200 1952 13252
rect 2004 13240 2010 13252
rect 2056 13240 2084 13271
rect 2222 13268 2228 13320
rect 2280 13268 2286 13320
rect 3234 13268 3240 13320
rect 3292 13268 3298 13320
rect 3329 13311 3387 13317
rect 3329 13277 3341 13311
rect 3375 13277 3387 13311
rect 3329 13271 3387 13277
rect 2498 13240 2504 13252
rect 2004 13212 2084 13240
rect 2332 13212 2504 13240
rect 2004 13200 2010 13212
rect 1581 13175 1639 13181
rect 1581 13141 1593 13175
rect 1627 13172 1639 13175
rect 2332 13172 2360 13212
rect 2498 13200 2504 13212
rect 2556 13240 2562 13252
rect 3344 13240 3372 13271
rect 4154 13268 4160 13320
rect 4212 13308 4218 13320
rect 5276 13317 5304 13348
rect 5920 13320 5948 13348
rect 5077 13311 5135 13317
rect 5077 13308 5089 13311
rect 4212 13280 5089 13308
rect 4212 13268 4218 13280
rect 5077 13277 5089 13280
rect 5123 13277 5135 13311
rect 5077 13271 5135 13277
rect 5261 13311 5319 13317
rect 5261 13277 5273 13311
rect 5307 13277 5319 13311
rect 5261 13271 5319 13277
rect 5353 13311 5411 13317
rect 5353 13277 5365 13311
rect 5399 13308 5411 13311
rect 5534 13308 5540 13320
rect 5399 13280 5540 13308
rect 5399 13277 5411 13280
rect 5353 13271 5411 13277
rect 2556 13212 3372 13240
rect 5092 13240 5120 13271
rect 5534 13268 5540 13280
rect 5592 13308 5598 13320
rect 5813 13311 5871 13317
rect 5813 13308 5825 13311
rect 5592 13280 5825 13308
rect 5592 13268 5598 13280
rect 5813 13277 5825 13280
rect 5859 13277 5871 13311
rect 5813 13271 5871 13277
rect 5902 13268 5908 13320
rect 5960 13308 5966 13320
rect 6089 13311 6147 13317
rect 6089 13308 6101 13311
rect 5960 13280 6101 13308
rect 5960 13268 5966 13280
rect 6089 13277 6101 13280
rect 6135 13277 6147 13311
rect 6089 13271 6147 13277
rect 6472 13308 6500 13416
rect 7098 13404 7104 13456
rect 7156 13444 7162 13456
rect 7374 13444 7380 13456
rect 7156 13416 7380 13444
rect 7156 13404 7162 13416
rect 7374 13404 7380 13416
rect 7432 13404 7438 13456
rect 7576 13444 7604 13472
rect 7484 13416 7604 13444
rect 6733 13311 6791 13317
rect 6733 13308 6745 13311
rect 6472 13280 6745 13308
rect 5997 13243 6055 13249
rect 5997 13240 6009 13243
rect 5092 13212 6009 13240
rect 2556 13200 2562 13212
rect 5997 13209 6009 13212
rect 6043 13209 6055 13243
rect 5997 13203 6055 13209
rect 6472 13184 6500 13280
rect 6733 13277 6745 13280
rect 6779 13277 6791 13311
rect 6733 13271 6791 13277
rect 7190 13268 7196 13320
rect 7248 13308 7254 13320
rect 7484 13317 7512 13416
rect 11054 13404 11060 13456
rect 11112 13444 11118 13456
rect 11112 13416 11652 13444
rect 11112 13404 11118 13416
rect 10781 13379 10839 13385
rect 7576 13348 10180 13376
rect 7469 13311 7527 13317
rect 7248 13280 7420 13308
rect 7248 13268 7254 13280
rect 7392 13249 7420 13280
rect 7469 13277 7481 13311
rect 7515 13277 7527 13311
rect 7469 13271 7527 13277
rect 7377 13243 7435 13249
rect 7377 13209 7389 13243
rect 7423 13209 7435 13243
rect 7377 13203 7435 13209
rect 1627 13144 2360 13172
rect 1627 13141 1639 13144
rect 1581 13135 1639 13141
rect 2406 13132 2412 13184
rect 2464 13132 2470 13184
rect 4890 13132 4896 13184
rect 4948 13132 4954 13184
rect 6454 13132 6460 13184
rect 6512 13132 6518 13184
rect 6546 13132 6552 13184
rect 6604 13132 6610 13184
rect 7576 13181 7604 13348
rect 10152 13320 10180 13348
rect 10781 13345 10793 13379
rect 10827 13376 10839 13379
rect 10827 13348 11468 13376
rect 10827 13345 10839 13348
rect 10781 13339 10839 13345
rect 7650 13268 7656 13320
rect 7708 13268 7714 13320
rect 8386 13268 8392 13320
rect 8444 13308 8450 13320
rect 8941 13311 8999 13317
rect 8941 13308 8953 13311
rect 8444 13280 8953 13308
rect 8444 13268 8450 13280
rect 8941 13277 8953 13280
rect 8987 13277 8999 13311
rect 8941 13271 8999 13277
rect 10134 13268 10140 13320
rect 10192 13268 10198 13320
rect 10686 13268 10692 13320
rect 10744 13268 10750 13320
rect 10870 13268 10876 13320
rect 10928 13268 10934 13320
rect 11440 13317 11468 13348
rect 11624 13320 11652 13416
rect 11425 13311 11483 13317
rect 11425 13277 11437 13311
rect 11471 13308 11483 13311
rect 11514 13308 11520 13320
rect 11471 13280 11520 13308
rect 11471 13277 11483 13280
rect 11425 13271 11483 13277
rect 11514 13268 11520 13280
rect 11572 13268 11578 13320
rect 11606 13268 11612 13320
rect 11664 13268 11670 13320
rect 12360 13317 12388 13472
rect 12621 13447 12679 13453
rect 12621 13413 12633 13447
rect 12667 13444 12679 13447
rect 13004 13444 13032 13472
rect 12667 13416 13032 13444
rect 12667 13413 12679 13416
rect 12621 13407 12679 13413
rect 12529 13379 12587 13385
rect 12529 13345 12541 13379
rect 12575 13376 12587 13379
rect 12897 13379 12955 13385
rect 12897 13376 12909 13379
rect 12575 13348 12909 13376
rect 12575 13345 12587 13348
rect 12529 13339 12587 13345
rect 12897 13345 12909 13348
rect 12943 13345 12955 13379
rect 13004 13376 13032 13416
rect 13265 13379 13323 13385
rect 13265 13376 13277 13379
rect 13004 13348 13277 13376
rect 12897 13339 12955 13345
rect 13265 13345 13277 13348
rect 13311 13345 13323 13379
rect 13265 13339 13323 13345
rect 12345 13311 12403 13317
rect 12345 13277 12357 13311
rect 12391 13277 12403 13311
rect 12345 13271 12403 13277
rect 8205 13243 8263 13249
rect 8205 13209 8217 13243
rect 8251 13240 8263 13243
rect 8294 13240 8300 13252
rect 8251 13212 8300 13240
rect 8251 13209 8263 13212
rect 8205 13203 8263 13209
rect 8294 13200 8300 13212
rect 8352 13240 8358 13252
rect 9033 13243 9091 13249
rect 9033 13240 9045 13243
rect 8352 13212 9045 13240
rect 8352 13200 8358 13212
rect 9033 13209 9045 13212
rect 9079 13209 9091 13243
rect 9033 13203 9091 13209
rect 9217 13243 9275 13249
rect 9217 13209 9229 13243
rect 9263 13209 9275 13243
rect 9217 13203 9275 13209
rect 7177 13175 7235 13181
rect 7177 13141 7189 13175
rect 7223 13172 7235 13175
rect 7561 13175 7619 13181
rect 7561 13172 7573 13175
rect 7223 13144 7573 13172
rect 7223 13141 7235 13144
rect 7177 13135 7235 13141
rect 7561 13141 7573 13144
rect 7607 13141 7619 13175
rect 7561 13135 7619 13141
rect 8110 13132 8116 13184
rect 8168 13172 8174 13184
rect 8405 13175 8463 13181
rect 8405 13172 8417 13175
rect 8168 13144 8417 13172
rect 8168 13132 8174 13144
rect 8405 13141 8417 13144
rect 8451 13172 8463 13175
rect 9232 13172 9260 13203
rect 10318 13200 10324 13252
rect 10376 13200 10382 13252
rect 10505 13243 10563 13249
rect 10505 13209 10517 13243
rect 10551 13240 10563 13243
rect 10888 13240 10916 13268
rect 10551 13212 10916 13240
rect 10551 13209 10563 13212
rect 10505 13203 10563 13209
rect 8451 13144 9260 13172
rect 11517 13175 11575 13181
rect 8451 13141 8463 13144
rect 8405 13135 8463 13141
rect 11517 13141 11529 13175
rect 11563 13172 11575 13175
rect 12544 13172 12572 13339
rect 12710 13268 12716 13320
rect 12768 13308 12774 13320
rect 12805 13311 12863 13317
rect 12805 13308 12817 13311
rect 12768 13280 12817 13308
rect 12768 13268 12774 13280
rect 12805 13277 12817 13280
rect 12851 13277 12863 13311
rect 12805 13271 12863 13277
rect 13449 13311 13507 13317
rect 13449 13277 13461 13311
rect 13495 13277 13507 13311
rect 13449 13271 13507 13277
rect 13464 13240 13492 13271
rect 13906 13268 13912 13320
rect 13964 13308 13970 13320
rect 14277 13311 14335 13317
rect 14277 13308 14289 13311
rect 13964 13280 14289 13308
rect 13964 13268 13970 13280
rect 14277 13277 14289 13280
rect 14323 13277 14335 13311
rect 14553 13311 14611 13317
rect 14553 13308 14565 13311
rect 14277 13271 14335 13277
rect 14384 13280 14565 13308
rect 13188 13212 13492 13240
rect 13188 13181 13216 13212
rect 14384 13184 14412 13280
rect 14553 13277 14565 13280
rect 14599 13277 14611 13311
rect 14553 13271 14611 13277
rect 15746 13268 15752 13320
rect 15804 13268 15810 13320
rect 11563 13144 12572 13172
rect 13173 13175 13231 13181
rect 11563 13141 11575 13144
rect 11517 13135 11575 13141
rect 13173 13141 13185 13175
rect 13219 13141 13231 13175
rect 13173 13135 13231 13141
rect 13630 13132 13636 13184
rect 13688 13132 13694 13184
rect 14366 13132 14372 13184
rect 14424 13132 14430 13184
rect 14461 13175 14519 13181
rect 14461 13141 14473 13175
rect 14507 13172 14519 13175
rect 14826 13172 14832 13184
rect 14507 13144 14832 13172
rect 14507 13141 14519 13144
rect 14461 13135 14519 13141
rect 14826 13132 14832 13144
rect 14884 13132 14890 13184
rect 15930 13132 15936 13184
rect 15988 13132 15994 13184
rect 1104 13082 16376 13104
rect 1104 13030 3519 13082
rect 3571 13030 3583 13082
rect 3635 13030 3647 13082
rect 3699 13030 3711 13082
rect 3763 13030 3775 13082
rect 3827 13030 7337 13082
rect 7389 13030 7401 13082
rect 7453 13030 7465 13082
rect 7517 13030 7529 13082
rect 7581 13030 7593 13082
rect 7645 13030 11155 13082
rect 11207 13030 11219 13082
rect 11271 13030 11283 13082
rect 11335 13030 11347 13082
rect 11399 13030 11411 13082
rect 11463 13030 14973 13082
rect 15025 13030 15037 13082
rect 15089 13030 15101 13082
rect 15153 13030 15165 13082
rect 15217 13030 15229 13082
rect 15281 13030 16376 13082
rect 1104 13008 16376 13030
rect 2498 12928 2504 12980
rect 2556 12928 2562 12980
rect 2682 12928 2688 12980
rect 2740 12928 2746 12980
rect 3234 12928 3240 12980
rect 3292 12928 3298 12980
rect 4890 12928 4896 12980
rect 4948 12928 4954 12980
rect 4982 12928 4988 12980
rect 5040 12928 5046 12980
rect 5534 12928 5540 12980
rect 5592 12928 5598 12980
rect 5905 12971 5963 12977
rect 5905 12937 5917 12971
rect 5951 12968 5963 12971
rect 6546 12968 6552 12980
rect 5951 12940 6552 12968
rect 5951 12937 5963 12940
rect 5905 12931 5963 12937
rect 6546 12928 6552 12940
rect 6604 12928 6610 12980
rect 7653 12971 7711 12977
rect 7653 12937 7665 12971
rect 7699 12968 7711 12971
rect 8110 12968 8116 12980
rect 7699 12940 8116 12968
rect 7699 12937 7711 12940
rect 7653 12931 7711 12937
rect 8110 12928 8116 12940
rect 8168 12928 8174 12980
rect 8294 12928 8300 12980
rect 8352 12928 8358 12980
rect 8757 12971 8815 12977
rect 8757 12937 8769 12971
rect 8803 12968 8815 12971
rect 8846 12968 8852 12980
rect 8803 12940 8852 12968
rect 8803 12937 8815 12940
rect 8757 12931 8815 12937
rect 8846 12928 8852 12940
rect 8904 12928 8910 12980
rect 10134 12928 10140 12980
rect 10192 12928 10198 12980
rect 10321 12971 10379 12977
rect 10321 12937 10333 12971
rect 10367 12968 10379 12971
rect 10686 12968 10692 12980
rect 10367 12940 10692 12968
rect 10367 12937 10379 12940
rect 10321 12931 10379 12937
rect 10686 12928 10692 12940
rect 10744 12928 10750 12980
rect 11514 12928 11520 12980
rect 11572 12928 11578 12980
rect 15746 12928 15752 12980
rect 15804 12928 15810 12980
rect 1394 12792 1400 12844
rect 1452 12792 1458 12844
rect 2516 12841 2544 12928
rect 2225 12835 2283 12841
rect 2225 12801 2237 12835
rect 2271 12832 2283 12835
rect 2501 12835 2559 12841
rect 2501 12832 2513 12835
rect 2271 12804 2513 12832
rect 2271 12801 2283 12804
rect 2225 12795 2283 12801
rect 2501 12801 2513 12804
rect 2547 12801 2559 12835
rect 2501 12795 2559 12801
rect 2685 12835 2743 12841
rect 2685 12801 2697 12835
rect 2731 12832 2743 12835
rect 3252 12832 3280 12928
rect 4908 12900 4936 12928
rect 4632 12872 4936 12900
rect 4632 12841 4660 12872
rect 2731 12804 3280 12832
rect 4617 12835 4675 12841
rect 2731 12801 2743 12804
rect 2685 12795 2743 12801
rect 4617 12801 4629 12835
rect 4663 12801 4675 12835
rect 4617 12795 4675 12801
rect 4801 12835 4859 12841
rect 4801 12801 4813 12835
rect 4847 12832 4859 12835
rect 5000 12832 5028 12928
rect 7285 12903 7343 12909
rect 7285 12900 7297 12903
rect 6012 12872 7297 12900
rect 4847 12804 5028 12832
rect 4847 12801 4859 12804
rect 4801 12795 4859 12801
rect 5718 12792 5724 12844
rect 5776 12792 5782 12844
rect 6012 12841 6040 12872
rect 7285 12869 7297 12872
rect 7331 12900 7343 12903
rect 8389 12903 8447 12909
rect 8389 12900 8401 12903
rect 7331 12872 7512 12900
rect 7331 12869 7343 12872
rect 7285 12863 7343 12869
rect 7484 12844 7512 12872
rect 7576 12872 8156 12900
rect 5997 12835 6055 12841
rect 5997 12801 6009 12835
rect 6043 12801 6055 12835
rect 7193 12835 7251 12841
rect 7193 12832 7205 12835
rect 5997 12795 6055 12801
rect 6840 12804 7205 12832
rect 1854 12724 1860 12776
rect 1912 12764 1918 12776
rect 2038 12764 2044 12776
rect 1912 12736 2044 12764
rect 1912 12724 1918 12736
rect 2038 12724 2044 12736
rect 2096 12764 2102 12776
rect 2409 12767 2467 12773
rect 2409 12764 2421 12767
rect 2096 12736 2421 12764
rect 2096 12724 2102 12736
rect 2409 12733 2421 12736
rect 2455 12733 2467 12767
rect 2409 12727 2467 12733
rect 1581 12699 1639 12705
rect 1581 12665 1593 12699
rect 1627 12696 1639 12699
rect 6840 12696 6868 12804
rect 7193 12801 7205 12804
rect 7239 12801 7251 12835
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 7193 12795 7251 12801
rect 7300 12804 7389 12832
rect 6917 12767 6975 12773
rect 6917 12733 6929 12767
rect 6963 12764 6975 12767
rect 7098 12764 7104 12776
rect 6963 12736 7104 12764
rect 6963 12733 6975 12736
rect 6917 12727 6975 12733
rect 1627 12668 6868 12696
rect 1627 12665 1639 12668
rect 1581 12659 1639 12665
rect 1670 12588 1676 12640
rect 1728 12628 1734 12640
rect 2041 12631 2099 12637
rect 2041 12628 2053 12631
rect 1728 12600 2053 12628
rect 1728 12588 1734 12600
rect 2041 12597 2053 12600
rect 2087 12628 2099 12631
rect 2222 12628 2228 12640
rect 2087 12600 2228 12628
rect 2087 12597 2099 12600
rect 2041 12591 2099 12597
rect 2222 12588 2228 12600
rect 2280 12588 2286 12640
rect 4246 12588 4252 12640
rect 4304 12628 4310 12640
rect 4709 12631 4767 12637
rect 4709 12628 4721 12631
rect 4304 12600 4721 12628
rect 4304 12588 4310 12600
rect 4709 12597 4721 12600
rect 4755 12597 4767 12631
rect 4709 12591 4767 12597
rect 6546 12588 6552 12640
rect 6604 12628 6610 12640
rect 6932 12628 6960 12727
rect 7098 12724 7104 12736
rect 7156 12724 7162 12776
rect 7208 12696 7236 12795
rect 7300 12776 7328 12804
rect 7377 12801 7389 12804
rect 7423 12801 7435 12835
rect 7377 12795 7435 12801
rect 7466 12792 7472 12844
rect 7524 12792 7530 12844
rect 7282 12724 7288 12776
rect 7340 12724 7346 12776
rect 7576 12696 7604 12872
rect 7745 12835 7803 12841
rect 7745 12801 7757 12835
rect 7791 12801 7803 12835
rect 7745 12795 7803 12801
rect 7208 12668 7604 12696
rect 7760 12696 7788 12795
rect 7834 12792 7840 12844
rect 7892 12792 7898 12844
rect 7926 12792 7932 12844
rect 7984 12792 7990 12844
rect 8128 12841 8156 12872
rect 8312 12872 8401 12900
rect 8312 12844 8340 12872
rect 8389 12869 8401 12872
rect 8435 12869 8447 12903
rect 8389 12863 8447 12869
rect 8605 12903 8663 12909
rect 8605 12869 8617 12903
rect 8651 12900 8663 12903
rect 9122 12900 9128 12912
rect 8651 12872 9128 12900
rect 8651 12869 8663 12872
rect 8605 12863 8663 12869
rect 9122 12860 9128 12872
rect 9180 12860 9186 12912
rect 8021 12835 8079 12841
rect 8021 12801 8033 12835
rect 8067 12801 8079 12835
rect 8021 12795 8079 12801
rect 8113 12835 8171 12841
rect 8113 12801 8125 12835
rect 8159 12801 8171 12835
rect 8113 12795 8171 12801
rect 7852 12764 7880 12792
rect 8036 12764 8064 12795
rect 7852 12736 8064 12764
rect 8128 12764 8156 12795
rect 8294 12792 8300 12844
rect 8352 12792 8358 12844
rect 10152 12841 10180 12928
rect 10137 12835 10195 12841
rect 10137 12801 10149 12835
rect 10183 12801 10195 12835
rect 10137 12795 10195 12801
rect 10318 12792 10324 12844
rect 10376 12792 10382 12844
rect 11532 12832 11560 12928
rect 11701 12835 11759 12841
rect 11701 12832 11713 12835
rect 11532 12804 11713 12832
rect 11701 12801 11713 12804
rect 11747 12801 11759 12835
rect 11701 12795 11759 12801
rect 13449 12835 13507 12841
rect 13449 12801 13461 12835
rect 13495 12832 13507 12835
rect 13630 12832 13636 12844
rect 13495 12804 13636 12832
rect 13495 12801 13507 12804
rect 13449 12795 13507 12801
rect 13630 12792 13636 12804
rect 13688 12792 13694 12844
rect 14553 12835 14611 12841
rect 14553 12801 14565 12835
rect 14599 12832 14611 12835
rect 14826 12832 14832 12844
rect 14599 12804 14832 12832
rect 14599 12801 14611 12804
rect 14553 12795 14611 12801
rect 14826 12792 14832 12804
rect 14884 12792 14890 12844
rect 8128 12736 8616 12764
rect 8294 12696 8300 12708
rect 7760 12668 8300 12696
rect 8294 12656 8300 12668
rect 8352 12656 8358 12708
rect 8588 12640 8616 12736
rect 10042 12724 10048 12776
rect 10100 12764 10106 12776
rect 10336 12764 10364 12792
rect 10100 12736 10364 12764
rect 10100 12724 10106 12736
rect 11606 12724 11612 12776
rect 11664 12724 11670 12776
rect 13354 12724 13360 12776
rect 13412 12724 13418 12776
rect 14366 12764 14372 12776
rect 13832 12736 14372 12764
rect 13832 12705 13860 12736
rect 14366 12724 14372 12736
rect 14424 12764 14430 12776
rect 14461 12767 14519 12773
rect 14461 12764 14473 12767
rect 14424 12736 14473 12764
rect 14424 12724 14430 12736
rect 14461 12733 14473 12736
rect 14507 12733 14519 12767
rect 14461 12727 14519 12733
rect 14921 12767 14979 12773
rect 14921 12733 14933 12767
rect 14967 12764 14979 12767
rect 15764 12764 15792 12928
rect 14967 12736 15792 12764
rect 14967 12733 14979 12736
rect 14921 12727 14979 12733
rect 13817 12699 13875 12705
rect 13817 12665 13829 12699
rect 13863 12665 13875 12699
rect 13817 12659 13875 12665
rect 6604 12600 6960 12628
rect 7009 12631 7067 12637
rect 6604 12588 6610 12600
rect 7009 12597 7021 12631
rect 7055 12628 7067 12631
rect 7834 12628 7840 12640
rect 7055 12600 7840 12628
rect 7055 12597 7067 12600
rect 7009 12591 7067 12597
rect 7834 12588 7840 12600
rect 7892 12588 7898 12640
rect 8570 12588 8576 12640
rect 8628 12588 8634 12640
rect 12066 12588 12072 12640
rect 12124 12588 12130 12640
rect 1104 12538 16376 12560
rect 1104 12486 2859 12538
rect 2911 12486 2923 12538
rect 2975 12486 2987 12538
rect 3039 12486 3051 12538
rect 3103 12486 3115 12538
rect 3167 12486 6677 12538
rect 6729 12486 6741 12538
rect 6793 12486 6805 12538
rect 6857 12486 6869 12538
rect 6921 12486 6933 12538
rect 6985 12486 10495 12538
rect 10547 12486 10559 12538
rect 10611 12486 10623 12538
rect 10675 12486 10687 12538
rect 10739 12486 10751 12538
rect 10803 12486 14313 12538
rect 14365 12486 14377 12538
rect 14429 12486 14441 12538
rect 14493 12486 14505 12538
rect 14557 12486 14569 12538
rect 14621 12486 16376 12538
rect 1104 12464 16376 12486
rect 2038 12384 2044 12436
rect 2096 12384 2102 12436
rect 4433 12427 4491 12433
rect 4433 12393 4445 12427
rect 4479 12424 4491 12427
rect 5074 12424 5080 12436
rect 4479 12396 5080 12424
rect 4479 12393 4491 12396
rect 4433 12387 4491 12393
rect 2225 12359 2283 12365
rect 2225 12325 2237 12359
rect 2271 12325 2283 12359
rect 2225 12319 2283 12325
rect 2240 12288 2268 12319
rect 4540 12297 4568 12396
rect 5074 12384 5080 12396
rect 5132 12384 5138 12436
rect 5718 12384 5724 12436
rect 5776 12384 5782 12436
rect 5902 12384 5908 12436
rect 5960 12384 5966 12436
rect 7929 12427 7987 12433
rect 7929 12424 7941 12427
rect 7116 12396 7941 12424
rect 5736 12356 5764 12384
rect 5644 12328 5764 12356
rect 5920 12356 5948 12384
rect 7116 12368 7144 12396
rect 7929 12393 7941 12396
rect 7975 12393 7987 12427
rect 7929 12387 7987 12393
rect 8297 12427 8355 12433
rect 8297 12393 8309 12427
rect 8343 12424 8355 12427
rect 8386 12424 8392 12436
rect 8343 12396 8392 12424
rect 8343 12393 8355 12396
rect 8297 12387 8355 12393
rect 8386 12384 8392 12396
rect 8444 12384 8450 12436
rect 9493 12427 9551 12433
rect 9493 12393 9505 12427
rect 9539 12424 9551 12427
rect 10042 12424 10048 12436
rect 9539 12396 10048 12424
rect 9539 12393 9551 12396
rect 9493 12387 9551 12393
rect 10042 12384 10048 12396
rect 10100 12384 10106 12436
rect 12342 12384 12348 12436
rect 12400 12424 12406 12436
rect 12400 12396 13032 12424
rect 12400 12384 12406 12396
rect 5920 12328 6408 12356
rect 2409 12291 2467 12297
rect 2409 12288 2421 12291
rect 2240 12260 2421 12288
rect 2409 12257 2421 12260
rect 2455 12257 2467 12291
rect 2409 12251 2467 12257
rect 2869 12291 2927 12297
rect 2869 12257 2881 12291
rect 2915 12257 2927 12291
rect 2869 12251 2927 12257
rect 4525 12291 4583 12297
rect 4525 12257 4537 12291
rect 4571 12257 4583 12291
rect 4525 12251 4583 12257
rect 5261 12291 5319 12297
rect 5261 12257 5273 12291
rect 5307 12257 5319 12291
rect 5261 12251 5319 12257
rect 1670 12180 1676 12232
rect 1728 12180 1734 12232
rect 2498 12180 2504 12232
rect 2556 12180 2562 12232
rect 2884 12220 2912 12251
rect 3418 12220 3424 12232
rect 2884 12192 3424 12220
rect 3418 12180 3424 12192
rect 3476 12180 3482 12232
rect 3973 12223 4031 12229
rect 3973 12189 3985 12223
rect 4019 12220 4031 12223
rect 4154 12220 4160 12232
rect 4019 12192 4160 12220
rect 4019 12189 4031 12192
rect 3973 12183 4031 12189
rect 4154 12180 4160 12192
rect 4212 12180 4218 12232
rect 4246 12180 4252 12232
rect 4304 12180 4310 12232
rect 4706 12180 4712 12232
rect 4764 12180 4770 12232
rect 1946 12112 1952 12164
rect 2004 12152 2010 12164
rect 2041 12155 2099 12161
rect 2041 12152 2053 12155
rect 2004 12124 2053 12152
rect 2004 12112 2010 12124
rect 2041 12121 2053 12124
rect 2087 12152 2099 12155
rect 2222 12152 2228 12164
rect 2087 12124 2228 12152
rect 2087 12121 2099 12124
rect 2041 12115 2099 12121
rect 2222 12112 2228 12124
rect 2280 12112 2286 12164
rect 3234 12112 3240 12164
rect 3292 12152 3298 12164
rect 5276 12152 5304 12251
rect 5644 12229 5672 12328
rect 5721 12291 5779 12297
rect 5721 12257 5733 12291
rect 5767 12288 5779 12291
rect 6273 12291 6331 12297
rect 6273 12288 6285 12291
rect 5767 12260 6285 12288
rect 5767 12257 5779 12260
rect 5721 12251 5779 12257
rect 6273 12257 6285 12260
rect 6319 12257 6331 12291
rect 6273 12251 6331 12257
rect 5629 12223 5687 12229
rect 5629 12189 5641 12223
rect 5675 12189 5687 12223
rect 5629 12183 5687 12189
rect 5902 12180 5908 12232
rect 5960 12180 5966 12232
rect 5994 12180 6000 12232
rect 6052 12220 6058 12232
rect 6089 12223 6147 12229
rect 6089 12220 6101 12223
rect 6052 12192 6101 12220
rect 6052 12180 6058 12192
rect 6089 12189 6101 12192
rect 6135 12189 6147 12223
rect 6089 12183 6147 12189
rect 3292 12124 5304 12152
rect 6104 12152 6132 12183
rect 6178 12180 6184 12232
rect 6236 12180 6242 12232
rect 6380 12229 6408 12328
rect 7098 12316 7104 12368
rect 7156 12316 7162 12368
rect 8018 12356 8024 12368
rect 7760 12328 8024 12356
rect 7760 12300 7788 12328
rect 8018 12316 8024 12328
rect 8076 12316 8082 12368
rect 11974 12316 11980 12368
rect 12032 12356 12038 12368
rect 12529 12359 12587 12365
rect 12529 12356 12541 12359
rect 12032 12328 12541 12356
rect 12032 12316 12038 12328
rect 12529 12325 12541 12328
rect 12575 12325 12587 12359
rect 12529 12319 12587 12325
rect 7742 12248 7748 12300
rect 7800 12248 7806 12300
rect 9030 12248 9036 12300
rect 9088 12248 9094 12300
rect 6365 12223 6423 12229
rect 6365 12189 6377 12223
rect 6411 12189 6423 12223
rect 6365 12183 6423 12189
rect 7466 12180 7472 12232
rect 7524 12220 7530 12232
rect 7653 12223 7711 12229
rect 7653 12220 7665 12223
rect 7524 12192 7665 12220
rect 7524 12180 7530 12192
rect 7653 12189 7665 12192
rect 7699 12220 7711 12223
rect 7760 12220 7788 12248
rect 7699 12192 7788 12220
rect 7699 12189 7711 12192
rect 7653 12183 7711 12189
rect 7834 12180 7840 12232
rect 7892 12180 7898 12232
rect 7929 12223 7987 12229
rect 7929 12189 7941 12223
rect 7975 12189 7987 12223
rect 7929 12183 7987 12189
rect 6546 12152 6552 12164
rect 6104 12124 6552 12152
rect 3292 12112 3298 12124
rect 6546 12112 6552 12124
rect 6604 12112 6610 12164
rect 7745 12155 7803 12161
rect 7745 12121 7757 12155
rect 7791 12152 7803 12155
rect 7944 12152 7972 12183
rect 8018 12180 8024 12232
rect 8076 12180 8082 12232
rect 9122 12180 9128 12232
rect 9180 12180 9186 12232
rect 11885 12223 11943 12229
rect 11885 12220 11897 12223
rect 10888 12192 11897 12220
rect 9140 12152 9168 12180
rect 7791 12124 9168 12152
rect 7791 12121 7803 12124
rect 7745 12115 7803 12121
rect 10888 12096 10916 12192
rect 11885 12189 11897 12192
rect 11931 12189 11943 12223
rect 11885 12183 11943 12189
rect 11900 12152 11928 12183
rect 12066 12180 12072 12232
rect 12124 12220 12130 12232
rect 13004 12229 13032 12396
rect 13906 12384 13912 12436
rect 13964 12384 13970 12436
rect 13630 12316 13636 12368
rect 13688 12356 13694 12368
rect 13725 12359 13783 12365
rect 13725 12356 13737 12359
rect 13688 12328 13737 12356
rect 13688 12316 13694 12328
rect 13725 12325 13737 12328
rect 13771 12325 13783 12359
rect 13725 12319 13783 12325
rect 12161 12223 12219 12229
rect 12161 12220 12173 12223
rect 12124 12192 12173 12220
rect 12124 12180 12130 12192
rect 12161 12189 12173 12192
rect 12207 12220 12219 12223
rect 12437 12223 12495 12229
rect 12437 12220 12449 12223
rect 12207 12192 12449 12220
rect 12207 12189 12219 12192
rect 12161 12183 12219 12189
rect 12437 12189 12449 12192
rect 12483 12189 12495 12223
rect 12437 12183 12495 12189
rect 12805 12223 12863 12229
rect 12805 12189 12817 12223
rect 12851 12189 12863 12223
rect 12805 12183 12863 12189
rect 12989 12223 13047 12229
rect 12989 12189 13001 12223
rect 13035 12189 13047 12223
rect 12989 12183 13047 12189
rect 12713 12155 12771 12161
rect 12713 12152 12725 12155
rect 11900 12124 12725 12152
rect 12713 12121 12725 12124
rect 12759 12121 12771 12155
rect 12713 12115 12771 12121
rect 3605 12087 3663 12093
rect 3605 12053 3617 12087
rect 3651 12084 3663 12087
rect 4062 12084 4068 12096
rect 3651 12056 4068 12084
rect 3651 12053 3663 12056
rect 3605 12047 3663 12053
rect 4062 12044 4068 12056
rect 4120 12044 4126 12096
rect 4893 12087 4951 12093
rect 4893 12053 4905 12087
rect 4939 12084 4951 12087
rect 9950 12084 9956 12096
rect 4939 12056 9956 12084
rect 4939 12053 4951 12056
rect 4893 12047 4951 12053
rect 9950 12044 9956 12056
rect 10008 12044 10014 12096
rect 10870 12044 10876 12096
rect 10928 12044 10934 12096
rect 12437 12087 12495 12093
rect 12437 12053 12449 12087
rect 12483 12084 12495 12087
rect 12820 12084 12848 12183
rect 13446 12112 13452 12164
rect 13504 12112 13510 12164
rect 12483 12056 12848 12084
rect 12483 12053 12495 12056
rect 12437 12047 12495 12053
rect 12894 12044 12900 12096
rect 12952 12044 12958 12096
rect 1104 11994 16376 12016
rect 1104 11942 3519 11994
rect 3571 11942 3583 11994
rect 3635 11942 3647 11994
rect 3699 11942 3711 11994
rect 3763 11942 3775 11994
rect 3827 11942 7337 11994
rect 7389 11942 7401 11994
rect 7453 11942 7465 11994
rect 7517 11942 7529 11994
rect 7581 11942 7593 11994
rect 7645 11942 11155 11994
rect 11207 11942 11219 11994
rect 11271 11942 11283 11994
rect 11335 11942 11347 11994
rect 11399 11942 11411 11994
rect 11463 11942 14973 11994
rect 15025 11942 15037 11994
rect 15089 11942 15101 11994
rect 15153 11942 15165 11994
rect 15217 11942 15229 11994
rect 15281 11942 16376 11994
rect 1104 11920 16376 11942
rect 3234 11840 3240 11892
rect 3292 11840 3298 11892
rect 3418 11840 3424 11892
rect 3476 11840 3482 11892
rect 4062 11840 4068 11892
rect 4120 11840 4126 11892
rect 4157 11883 4215 11889
rect 4157 11849 4169 11883
rect 4203 11880 4215 11883
rect 4706 11880 4712 11892
rect 4203 11852 4712 11880
rect 4203 11849 4215 11852
rect 4157 11843 4215 11849
rect 4706 11840 4712 11852
rect 4764 11840 4770 11892
rect 8757 11883 8815 11889
rect 8404 11852 8708 11880
rect 3252 11753 3280 11840
rect 3436 11753 3464 11840
rect 4080 11753 4108 11840
rect 4246 11772 4252 11824
rect 4304 11812 4310 11824
rect 4341 11815 4399 11821
rect 4341 11812 4353 11815
rect 4304 11784 4353 11812
rect 4304 11772 4310 11784
rect 4341 11781 4353 11784
rect 4387 11781 4399 11815
rect 4341 11775 4399 11781
rect 7190 11772 7196 11824
rect 7248 11812 7254 11824
rect 7558 11812 7564 11824
rect 7248 11784 7564 11812
rect 7248 11772 7254 11784
rect 7558 11772 7564 11784
rect 7616 11812 7622 11824
rect 8404 11821 8432 11852
rect 8389 11815 8447 11821
rect 8389 11812 8401 11815
rect 7616 11784 8401 11812
rect 7616 11772 7622 11784
rect 8389 11781 8401 11784
rect 8435 11781 8447 11815
rect 8589 11815 8647 11821
rect 8589 11812 8601 11815
rect 8389 11775 8447 11781
rect 8496 11784 8601 11812
rect 3237 11747 3295 11753
rect 3237 11713 3249 11747
rect 3283 11713 3295 11747
rect 3237 11707 3295 11713
rect 3421 11747 3479 11753
rect 3421 11713 3433 11747
rect 3467 11713 3479 11747
rect 3421 11707 3479 11713
rect 3697 11747 3755 11753
rect 3697 11713 3709 11747
rect 3743 11744 3755 11747
rect 4065 11747 4123 11753
rect 4065 11744 4077 11747
rect 3743 11716 4077 11744
rect 3743 11713 3755 11716
rect 3697 11707 3755 11713
rect 4065 11713 4077 11716
rect 4111 11713 4123 11747
rect 4065 11707 4123 11713
rect 4154 11704 4160 11756
rect 4212 11704 4218 11756
rect 8496 11688 8524 11784
rect 8589 11781 8601 11784
rect 8635 11781 8647 11815
rect 8680 11812 8708 11852
rect 8757 11849 8769 11883
rect 8803 11880 8815 11883
rect 9030 11880 9036 11892
rect 8803 11852 9036 11880
rect 8803 11849 8815 11852
rect 8757 11843 8815 11849
rect 9030 11840 9036 11852
rect 9088 11840 9094 11892
rect 10705 11883 10763 11889
rect 10705 11880 10717 11883
rect 10152 11852 10717 11880
rect 8846 11812 8852 11824
rect 8680 11784 8852 11812
rect 8589 11775 8647 11781
rect 8846 11772 8852 11784
rect 8904 11772 8910 11824
rect 9677 11815 9735 11821
rect 9677 11781 9689 11815
rect 9723 11812 9735 11815
rect 9723 11784 10088 11812
rect 9723 11781 9735 11784
rect 9677 11775 9735 11781
rect 9585 11747 9643 11753
rect 9585 11744 9597 11747
rect 8680 11716 9597 11744
rect 3329 11679 3387 11685
rect 3329 11645 3341 11679
rect 3375 11676 3387 11679
rect 3513 11679 3571 11685
rect 3513 11676 3525 11679
rect 3375 11648 3525 11676
rect 3375 11645 3387 11648
rect 3329 11639 3387 11645
rect 3513 11645 3525 11648
rect 3559 11645 3571 11679
rect 3513 11639 3571 11645
rect 8478 11636 8484 11688
rect 8536 11636 8542 11688
rect 8680 11552 8708 11716
rect 9585 11713 9597 11716
rect 9631 11713 9643 11747
rect 9769 11747 9827 11753
rect 9769 11744 9781 11747
rect 9585 11707 9643 11713
rect 9692 11716 9781 11744
rect 3878 11500 3884 11552
rect 3936 11500 3942 11552
rect 6638 11500 6644 11552
rect 6696 11540 6702 11552
rect 7466 11540 7472 11552
rect 6696 11512 7472 11540
rect 6696 11500 6702 11512
rect 7466 11500 7472 11512
rect 7524 11500 7530 11552
rect 7650 11500 7656 11552
rect 7708 11540 7714 11552
rect 8570 11540 8576 11552
rect 7708 11512 8576 11540
rect 7708 11500 7714 11512
rect 8570 11500 8576 11512
rect 8628 11500 8634 11552
rect 8662 11500 8668 11552
rect 8720 11500 8726 11552
rect 9600 11540 9628 11707
rect 9692 11620 9720 11716
rect 9769 11713 9781 11716
rect 9815 11713 9827 11747
rect 9769 11707 9827 11713
rect 9950 11704 9956 11756
rect 10008 11704 10014 11756
rect 10060 11753 10088 11784
rect 10045 11747 10103 11753
rect 10045 11713 10057 11747
rect 10091 11713 10103 11747
rect 10045 11707 10103 11713
rect 9968 11676 9996 11704
rect 10152 11685 10180 11852
rect 10705 11849 10717 11852
rect 10751 11849 10763 11883
rect 10705 11843 10763 11849
rect 10870 11840 10876 11892
rect 10928 11840 10934 11892
rect 11609 11883 11667 11889
rect 11609 11849 11621 11883
rect 11655 11880 11667 11883
rect 11974 11880 11980 11892
rect 11655 11852 11980 11880
rect 11655 11849 11667 11852
rect 11609 11843 11667 11849
rect 11974 11840 11980 11852
rect 12032 11880 12038 11892
rect 12250 11880 12256 11892
rect 12032 11852 12256 11880
rect 12032 11840 12038 11852
rect 12250 11840 12256 11852
rect 12308 11840 12314 11892
rect 12894 11840 12900 11892
rect 12952 11840 12958 11892
rect 14826 11840 14832 11892
rect 14884 11840 14890 11892
rect 10505 11815 10563 11821
rect 10505 11812 10517 11815
rect 10244 11784 10517 11812
rect 10137 11679 10195 11685
rect 10137 11676 10149 11679
rect 9968 11648 10149 11676
rect 10137 11645 10149 11648
rect 10183 11645 10195 11679
rect 10137 11639 10195 11645
rect 9674 11568 9680 11620
rect 9732 11608 9738 11620
rect 10244 11608 10272 11784
rect 10505 11781 10517 11784
rect 10551 11781 10563 11815
rect 10505 11775 10563 11781
rect 11514 11744 11520 11756
rect 10428 11716 11520 11744
rect 10428 11685 10456 11716
rect 11514 11704 11520 11716
rect 11572 11704 11578 11756
rect 11698 11704 11704 11756
rect 11756 11704 11762 11756
rect 12912 11744 12940 11840
rect 15197 11815 15255 11821
rect 15197 11812 15209 11815
rect 14844 11784 15209 11812
rect 14844 11756 14872 11784
rect 15197 11781 15209 11784
rect 15243 11781 15255 11815
rect 15197 11775 15255 11781
rect 14090 11744 14096 11756
rect 12912 11716 14096 11744
rect 14090 11704 14096 11716
rect 14148 11744 14154 11756
rect 14369 11747 14427 11753
rect 14369 11744 14381 11747
rect 14148 11716 14381 11744
rect 14148 11704 14154 11716
rect 14369 11713 14381 11716
rect 14415 11713 14427 11747
rect 14369 11707 14427 11713
rect 14826 11704 14832 11756
rect 14884 11704 14890 11756
rect 15010 11704 15016 11756
rect 15068 11704 15074 11756
rect 15289 11747 15347 11753
rect 15289 11713 15301 11747
rect 15335 11713 15347 11747
rect 15289 11707 15347 11713
rect 10413 11679 10471 11685
rect 10413 11645 10425 11679
rect 10459 11645 10471 11679
rect 14277 11679 14335 11685
rect 14277 11676 14289 11679
rect 10413 11639 10471 11645
rect 14200 11648 14289 11676
rect 9732 11580 10272 11608
rect 9732 11568 9738 11580
rect 14200 11552 14228 11648
rect 14277 11645 14289 11648
rect 14323 11645 14335 11679
rect 14277 11639 14335 11645
rect 14737 11679 14795 11685
rect 14737 11645 14749 11679
rect 14783 11676 14795 11679
rect 15194 11676 15200 11688
rect 14783 11648 15200 11676
rect 14783 11645 14795 11648
rect 14737 11639 14795 11645
rect 15194 11636 15200 11648
rect 15252 11676 15258 11688
rect 15304 11676 15332 11707
rect 15252 11648 15332 11676
rect 15252 11636 15258 11648
rect 10689 11543 10747 11549
rect 10689 11540 10701 11543
rect 9600 11512 10701 11540
rect 10689 11509 10701 11512
rect 10735 11509 10747 11543
rect 10689 11503 10747 11509
rect 14182 11500 14188 11552
rect 14240 11500 14246 11552
rect 1104 11450 16376 11472
rect 1104 11398 2859 11450
rect 2911 11398 2923 11450
rect 2975 11398 2987 11450
rect 3039 11398 3051 11450
rect 3103 11398 3115 11450
rect 3167 11398 6677 11450
rect 6729 11398 6741 11450
rect 6793 11398 6805 11450
rect 6857 11398 6869 11450
rect 6921 11398 6933 11450
rect 6985 11398 10495 11450
rect 10547 11398 10559 11450
rect 10611 11398 10623 11450
rect 10675 11398 10687 11450
rect 10739 11398 10751 11450
rect 10803 11398 14313 11450
rect 14365 11398 14377 11450
rect 14429 11398 14441 11450
rect 14493 11398 14505 11450
rect 14557 11398 14569 11450
rect 14621 11398 16376 11450
rect 1104 11376 16376 11398
rect 6454 11296 6460 11348
rect 6512 11296 6518 11348
rect 7098 11296 7104 11348
rect 7156 11336 7162 11348
rect 8297 11339 8355 11345
rect 8297 11336 8309 11339
rect 7156 11308 8309 11336
rect 7156 11296 7162 11308
rect 8297 11305 8309 11308
rect 8343 11305 8355 11339
rect 8297 11299 8355 11305
rect 8662 11296 8668 11348
rect 8720 11296 8726 11348
rect 11793 11339 11851 11345
rect 11793 11305 11805 11339
rect 11839 11336 11851 11339
rect 14737 11339 14795 11345
rect 11839 11308 12204 11336
rect 11839 11305 11851 11308
rect 11793 11299 11851 11305
rect 1581 11271 1639 11277
rect 1581 11237 1593 11271
rect 1627 11268 1639 11271
rect 5810 11268 5816 11280
rect 1627 11240 5816 11268
rect 1627 11237 1639 11240
rect 1581 11231 1639 11237
rect 5810 11228 5816 11240
rect 5868 11228 5874 11280
rect 7742 11268 7748 11280
rect 7300 11240 7748 11268
rect 6730 11160 6736 11212
rect 6788 11200 6794 11212
rect 6788 11172 7052 11200
rect 6788 11160 6794 11172
rect 1394 11092 1400 11144
rect 1452 11092 1458 11144
rect 7024 11141 7052 11172
rect 7300 11141 7328 11240
rect 7742 11228 7748 11240
rect 7800 11228 7806 11280
rect 8113 11271 8171 11277
rect 8113 11237 8125 11271
rect 8159 11268 8171 11271
rect 9674 11268 9680 11280
rect 8159 11240 9680 11268
rect 8159 11237 8171 11240
rect 8113 11231 8171 11237
rect 9674 11228 9680 11240
rect 9732 11228 9738 11280
rect 11698 11268 11704 11280
rect 11440 11240 11704 11268
rect 11440 11209 11468 11240
rect 11698 11228 11704 11240
rect 11756 11268 11762 11280
rect 11756 11240 12112 11268
rect 11756 11228 11762 11240
rect 7377 11203 7435 11209
rect 7377 11169 7389 11203
rect 7423 11200 7435 11203
rect 8389 11203 8447 11209
rect 7423 11172 8248 11200
rect 7423 11169 7435 11172
rect 7377 11163 7435 11169
rect 6641 11135 6699 11141
rect 6641 11132 6653 11135
rect 6196 11104 6653 11132
rect 6196 11008 6224 11104
rect 6641 11101 6653 11104
rect 6687 11132 6699 11135
rect 6917 11135 6975 11141
rect 6917 11132 6929 11135
rect 6687 11104 6929 11132
rect 6687 11101 6699 11104
rect 6641 11095 6699 11101
rect 6917 11101 6929 11104
rect 6963 11101 6975 11135
rect 6917 11095 6975 11101
rect 7009 11135 7067 11141
rect 7009 11101 7021 11135
rect 7055 11132 7067 11135
rect 7285 11135 7343 11141
rect 7055 11104 7220 11132
rect 7055 11101 7067 11104
rect 7009 11095 7067 11101
rect 7098 11064 7104 11076
rect 6288 11036 7104 11064
rect 6288 11008 6316 11036
rect 7098 11024 7104 11036
rect 7156 11024 7162 11076
rect 7192 11064 7220 11104
rect 7285 11101 7297 11135
rect 7331 11101 7343 11135
rect 7285 11095 7343 11101
rect 7466 11092 7472 11144
rect 7524 11092 7530 11144
rect 7558 11092 7564 11144
rect 7616 11092 7622 11144
rect 7650 11092 7656 11144
rect 7708 11132 7714 11144
rect 7953 11135 8011 11141
rect 7953 11134 7965 11135
rect 7852 11132 7965 11134
rect 7708 11106 7965 11132
rect 7708 11104 7880 11106
rect 7944 11104 7965 11106
rect 7708 11092 7714 11104
rect 7953 11101 7965 11104
rect 7999 11101 8011 11135
rect 8220 11134 8248 11172
rect 8389 11169 8401 11203
rect 8435 11200 8447 11203
rect 9033 11203 9091 11209
rect 9033 11200 9045 11203
rect 8435 11172 9045 11200
rect 8435 11169 8447 11172
rect 8389 11163 8447 11169
rect 9033 11169 9045 11172
rect 9079 11169 9091 11203
rect 9033 11163 9091 11169
rect 10965 11203 11023 11209
rect 10965 11169 10977 11203
rect 11011 11200 11023 11203
rect 11425 11203 11483 11209
rect 11425 11200 11437 11203
rect 11011 11172 11437 11200
rect 11011 11169 11023 11172
rect 10965 11163 11023 11169
rect 11425 11169 11437 11172
rect 11471 11169 11483 11203
rect 11425 11163 11483 11169
rect 8297 11135 8355 11141
rect 8297 11134 8309 11135
rect 8220 11106 8309 11134
rect 7953 11095 8011 11101
rect 8297 11101 8309 11106
rect 8343 11134 8355 11135
rect 8343 11132 8432 11134
rect 8478 11132 8484 11144
rect 8343 11106 8484 11132
rect 8343 11101 8355 11106
rect 8404 11104 8484 11106
rect 8297 11095 8355 11101
rect 8478 11092 8484 11104
rect 8536 11092 8542 11144
rect 8846 11092 8852 11144
rect 8904 11132 8910 11144
rect 8941 11135 8999 11141
rect 8941 11132 8953 11135
rect 8904 11104 8953 11132
rect 8904 11092 8910 11104
rect 8941 11101 8953 11104
rect 8987 11101 8999 11135
rect 11057 11135 11115 11141
rect 11057 11132 11069 11135
rect 8941 11095 8999 11101
rect 10612 11104 11069 11132
rect 7668 11064 7696 11092
rect 7192 11036 7696 11064
rect 7742 11024 7748 11076
rect 7800 11024 7806 11076
rect 7837 11067 7895 11073
rect 7837 11033 7849 11067
rect 7883 11033 7895 11067
rect 8496 11064 8524 11092
rect 10612 11073 10640 11104
rect 11057 11101 11069 11104
rect 11103 11101 11115 11135
rect 11241 11135 11299 11141
rect 11241 11132 11253 11135
rect 11057 11095 11115 11101
rect 11164 11104 11253 11132
rect 10597 11067 10655 11073
rect 10597 11064 10609 11067
rect 8496 11036 10609 11064
rect 7837 11027 7895 11033
rect 10597 11033 10609 11036
rect 10643 11033 10655 11067
rect 10597 11027 10655 11033
rect 10781 11067 10839 11073
rect 10781 11033 10793 11067
rect 10827 11064 10839 11067
rect 11164 11064 11192 11104
rect 11241 11101 11253 11104
rect 11287 11101 11299 11135
rect 11241 11095 11299 11101
rect 11514 11092 11520 11144
rect 11572 11132 11578 11144
rect 12084 11141 12112 11240
rect 12176 11141 12204 11308
rect 14737 11305 14749 11339
rect 14783 11336 14795 11339
rect 15010 11336 15016 11348
rect 14783 11308 15016 11336
rect 14783 11305 14795 11308
rect 14737 11299 14795 11305
rect 15010 11296 15016 11308
rect 15068 11296 15074 11348
rect 15194 11296 15200 11348
rect 15252 11296 15258 11348
rect 13814 11268 13820 11280
rect 12452 11240 13820 11268
rect 11609 11135 11667 11141
rect 11609 11132 11621 11135
rect 11572 11104 11621 11132
rect 11572 11092 11578 11104
rect 11609 11101 11621 11104
rect 11655 11101 11667 11135
rect 12069 11135 12127 11141
rect 11885 11126 11943 11131
rect 11609 11095 11667 11101
rect 11808 11125 11943 11126
rect 11808 11098 11897 11125
rect 11808 11064 11836 11098
rect 11885 11091 11897 11098
rect 11931 11091 11943 11125
rect 12069 11101 12081 11135
rect 12115 11101 12127 11135
rect 12069 11095 12127 11101
rect 12161 11135 12219 11141
rect 12161 11101 12173 11135
rect 12207 11101 12219 11135
rect 12161 11095 12219 11101
rect 12250 11092 12256 11144
rect 12308 11132 12314 11144
rect 12345 11135 12403 11141
rect 12345 11132 12357 11135
rect 12308 11104 12357 11132
rect 12308 11092 12314 11104
rect 12345 11101 12357 11104
rect 12391 11101 12403 11135
rect 12345 11095 12403 11101
rect 11885 11085 11943 11091
rect 12452 11064 12480 11240
rect 13814 11228 13820 11240
rect 13872 11228 13878 11280
rect 13449 11203 13507 11209
rect 13449 11169 13461 11203
rect 13495 11200 13507 11203
rect 13538 11200 13544 11212
rect 13495 11172 13544 11200
rect 13495 11169 13507 11172
rect 13449 11163 13507 11169
rect 13538 11160 13544 11172
rect 13596 11160 13602 11212
rect 13725 11203 13783 11209
rect 13725 11169 13737 11203
rect 13771 11200 13783 11203
rect 14182 11200 14188 11212
rect 13771 11172 14188 11200
rect 13771 11169 13783 11172
rect 13725 11163 13783 11169
rect 14182 11160 14188 11172
rect 14240 11200 14246 11212
rect 15212 11209 15240 11296
rect 15197 11203 15255 11209
rect 14240 11172 14596 11200
rect 14240 11160 14246 11172
rect 13354 11092 13360 11144
rect 13412 11092 13418 11144
rect 14090 11092 14096 11144
rect 14148 11132 14154 11144
rect 14568 11141 14596 11172
rect 15197 11169 15209 11203
rect 15243 11169 15255 11203
rect 15197 11163 15255 11169
rect 15654 11160 15660 11212
rect 15712 11160 15718 11212
rect 14369 11135 14427 11141
rect 14369 11132 14381 11135
rect 14148 11104 14381 11132
rect 14148 11092 14154 11104
rect 14369 11101 14381 11104
rect 14415 11101 14427 11135
rect 14369 11095 14427 11101
rect 14553 11135 14611 11141
rect 14553 11101 14565 11135
rect 14599 11101 14611 11135
rect 14553 11095 14611 11101
rect 14826 11092 14832 11144
rect 14884 11132 14890 11144
rect 15289 11135 15347 11141
rect 15289 11132 15301 11135
rect 14884 11104 15301 11132
rect 14884 11092 14890 11104
rect 15289 11101 15301 11104
rect 15335 11101 15347 11135
rect 15289 11095 15347 11101
rect 10827 11036 11192 11064
rect 11256 11036 11836 11064
rect 12268 11036 12480 11064
rect 12529 11067 12587 11073
rect 10827 11033 10839 11036
rect 10781 11027 10839 11033
rect 6178 10956 6184 11008
rect 6236 10956 6242 11008
rect 6270 10956 6276 11008
rect 6328 10956 6334 11008
rect 6454 10956 6460 11008
rect 6512 10996 6518 11008
rect 6733 10999 6791 11005
rect 6733 10996 6745 10999
rect 6512 10968 6745 10996
rect 6512 10956 6518 10968
rect 6733 10965 6745 10968
rect 6779 10965 6791 10999
rect 6733 10959 6791 10965
rect 7466 10956 7472 11008
rect 7524 10996 7530 11008
rect 7852 10996 7880 11027
rect 7926 10996 7932 11008
rect 7524 10968 7932 10996
rect 7524 10956 7530 10968
rect 7926 10956 7932 10968
rect 7984 10956 7990 11008
rect 9674 10956 9680 11008
rect 9732 10996 9738 11008
rect 10796 10996 10824 11027
rect 11256 11005 11284 11036
rect 9732 10968 10824 10996
rect 11241 10999 11299 11005
rect 9732 10956 9738 10968
rect 11241 10965 11253 10999
rect 11287 10965 11299 10999
rect 11241 10959 11299 10965
rect 12069 10999 12127 11005
rect 12069 10965 12081 10999
rect 12115 10996 12127 10999
rect 12268 10996 12296 11036
rect 12529 11033 12541 11067
rect 12575 11064 12587 11067
rect 13998 11064 14004 11076
rect 12575 11036 14004 11064
rect 12575 11033 12587 11036
rect 12529 11027 12587 11033
rect 13998 11024 14004 11036
rect 14056 11024 14062 11076
rect 12115 10968 12296 10996
rect 12115 10965 12127 10968
rect 12069 10959 12127 10965
rect 1104 10906 16376 10928
rect 1104 10854 3519 10906
rect 3571 10854 3583 10906
rect 3635 10854 3647 10906
rect 3699 10854 3711 10906
rect 3763 10854 3775 10906
rect 3827 10854 7337 10906
rect 7389 10854 7401 10906
rect 7453 10854 7465 10906
rect 7517 10854 7529 10906
rect 7581 10854 7593 10906
rect 7645 10854 11155 10906
rect 11207 10854 11219 10906
rect 11271 10854 11283 10906
rect 11335 10854 11347 10906
rect 11399 10854 11411 10906
rect 11463 10854 14973 10906
rect 15025 10854 15037 10906
rect 15089 10854 15101 10906
rect 15153 10854 15165 10906
rect 15217 10854 15229 10906
rect 15281 10854 16376 10906
rect 1104 10832 16376 10854
rect 3878 10752 3884 10804
rect 3936 10752 3942 10804
rect 4154 10752 4160 10804
rect 4212 10792 4218 10804
rect 5537 10795 5595 10801
rect 4212 10764 4568 10792
rect 4212 10752 4218 10764
rect 2406 10684 2412 10736
rect 2464 10724 2470 10736
rect 2501 10727 2559 10733
rect 2501 10724 2513 10727
rect 2464 10696 2513 10724
rect 2464 10684 2470 10696
rect 2501 10693 2513 10696
rect 2547 10693 2559 10727
rect 2501 10687 2559 10693
rect 3896 10724 3924 10752
rect 4540 10733 4568 10764
rect 5537 10761 5549 10795
rect 5583 10792 5595 10795
rect 5718 10792 5724 10804
rect 5583 10764 5724 10792
rect 5583 10761 5595 10764
rect 5537 10755 5595 10761
rect 5718 10752 5724 10764
rect 5776 10752 5782 10804
rect 6086 10752 6092 10804
rect 6144 10752 6150 10804
rect 9950 10752 9956 10804
rect 10008 10792 10014 10804
rect 13189 10795 13247 10801
rect 13189 10792 13201 10795
rect 10008 10764 13201 10792
rect 10008 10752 10014 10764
rect 13189 10761 13201 10764
rect 13235 10761 13247 10795
rect 13189 10755 13247 10761
rect 13357 10795 13415 10801
rect 13357 10761 13369 10795
rect 13403 10792 13415 10795
rect 13446 10792 13452 10804
rect 13403 10764 13452 10792
rect 13403 10761 13415 10764
rect 13357 10755 13415 10761
rect 13446 10752 13452 10764
rect 13504 10752 13510 10804
rect 15933 10795 15991 10801
rect 15933 10761 15945 10795
rect 15979 10792 15991 10795
rect 16022 10792 16028 10804
rect 15979 10764 16028 10792
rect 15979 10761 15991 10764
rect 15933 10755 15991 10761
rect 16022 10752 16028 10764
rect 16080 10752 16086 10804
rect 4433 10727 4491 10733
rect 4433 10724 4445 10727
rect 3896 10696 4445 10724
rect 934 10616 940 10668
rect 992 10656 998 10668
rect 1397 10659 1455 10665
rect 1397 10656 1409 10659
rect 992 10628 1409 10656
rect 992 10616 998 10628
rect 1397 10625 1409 10628
rect 1443 10625 1455 10659
rect 1397 10619 1455 10625
rect 2041 10659 2099 10665
rect 2041 10625 2053 10659
rect 2087 10656 2099 10659
rect 2424 10656 2452 10684
rect 2087 10628 2452 10656
rect 3697 10659 3755 10665
rect 2087 10625 2099 10628
rect 2041 10619 2099 10625
rect 3697 10625 3709 10659
rect 3743 10656 3755 10659
rect 3896 10656 3924 10696
rect 4433 10693 4445 10696
rect 4479 10693 4491 10727
rect 4433 10687 4491 10693
rect 4525 10727 4583 10733
rect 4525 10693 4537 10727
rect 4571 10724 4583 10727
rect 4614 10724 4620 10736
rect 4571 10696 4620 10724
rect 4571 10693 4583 10696
rect 4525 10687 4583 10693
rect 4614 10684 4620 10696
rect 4672 10684 4678 10736
rect 6104 10724 6132 10752
rect 6012 10696 6132 10724
rect 6012 10668 6040 10696
rect 6362 10684 6368 10736
rect 6420 10724 6426 10736
rect 12989 10727 13047 10733
rect 12989 10724 13001 10727
rect 6420 10696 7328 10724
rect 6420 10684 6426 10696
rect 3743 10628 3924 10656
rect 4801 10659 4859 10665
rect 3743 10625 3755 10628
rect 3697 10619 3755 10625
rect 4801 10625 4813 10659
rect 4847 10625 4859 10659
rect 4801 10619 4859 10625
rect 2133 10591 2191 10597
rect 2133 10557 2145 10591
rect 2179 10557 2191 10591
rect 2133 10551 2191 10557
rect 2148 10520 2176 10551
rect 2406 10548 2412 10600
rect 2464 10548 2470 10600
rect 2961 10591 3019 10597
rect 2961 10557 2973 10591
rect 3007 10588 3019 10591
rect 3789 10591 3847 10597
rect 3789 10588 3801 10591
rect 3007 10560 3801 10588
rect 3007 10557 3019 10560
rect 2961 10551 3019 10557
rect 3789 10557 3801 10560
rect 3835 10588 3847 10591
rect 4617 10591 4675 10597
rect 4617 10588 4629 10591
rect 3835 10560 4629 10588
rect 3835 10557 3847 10560
rect 3789 10551 3847 10557
rect 4617 10557 4629 10560
rect 4663 10557 4675 10591
rect 4617 10551 4675 10557
rect 2869 10523 2927 10529
rect 2869 10520 2881 10523
rect 2148 10492 2881 10520
rect 2869 10489 2881 10492
rect 2915 10520 2927 10523
rect 4430 10520 4436 10532
rect 2915 10492 3648 10520
rect 2915 10489 2927 10492
rect 2869 10483 2927 10489
rect 3620 10464 3648 10492
rect 3896 10492 4436 10520
rect 3896 10464 3924 10492
rect 4430 10480 4436 10492
rect 4488 10520 4494 10532
rect 4816 10520 4844 10619
rect 5074 10616 5080 10668
rect 5132 10656 5138 10668
rect 5353 10659 5411 10665
rect 5353 10656 5365 10659
rect 5132 10628 5365 10656
rect 5132 10616 5138 10628
rect 5353 10625 5365 10628
rect 5399 10656 5411 10659
rect 5629 10659 5687 10665
rect 5629 10656 5641 10659
rect 5399 10628 5641 10656
rect 5399 10625 5411 10628
rect 5353 10619 5411 10625
rect 5629 10625 5641 10628
rect 5675 10625 5687 10659
rect 5813 10659 5871 10665
rect 5813 10656 5825 10659
rect 5629 10619 5687 10625
rect 5736 10628 5825 10656
rect 5169 10591 5227 10597
rect 5169 10557 5181 10591
rect 5215 10588 5227 10591
rect 5215 10560 5672 10588
rect 5215 10557 5227 10560
rect 5169 10551 5227 10557
rect 4488 10492 4844 10520
rect 4488 10480 4494 10492
rect 5644 10464 5672 10560
rect 1581 10455 1639 10461
rect 1581 10421 1593 10455
rect 1627 10452 1639 10455
rect 3418 10452 3424 10464
rect 1627 10424 3424 10452
rect 1627 10421 1639 10424
rect 1581 10415 1639 10421
rect 3418 10412 3424 10424
rect 3476 10412 3482 10464
rect 3602 10412 3608 10464
rect 3660 10412 3666 10464
rect 3878 10412 3884 10464
rect 3936 10412 3942 10464
rect 4065 10455 4123 10461
rect 4065 10421 4077 10455
rect 4111 10452 4123 10455
rect 4338 10452 4344 10464
rect 4111 10424 4344 10452
rect 4111 10421 4123 10424
rect 4065 10415 4123 10421
rect 4338 10412 4344 10424
rect 4396 10412 4402 10464
rect 5626 10412 5632 10464
rect 5684 10412 5690 10464
rect 5736 10452 5764 10628
rect 5813 10625 5825 10628
rect 5859 10625 5871 10659
rect 5813 10619 5871 10625
rect 5994 10616 6000 10668
rect 6052 10616 6058 10668
rect 6086 10616 6092 10668
rect 6144 10616 6150 10668
rect 6546 10616 6552 10668
rect 6604 10656 6610 10668
rect 7300 10665 7328 10696
rect 12544 10696 13001 10724
rect 6641 10659 6699 10665
rect 6641 10656 6653 10659
rect 6604 10628 6653 10656
rect 6604 10616 6610 10628
rect 6641 10625 6653 10628
rect 6687 10625 6699 10659
rect 6641 10619 6699 10625
rect 7285 10659 7343 10665
rect 7285 10625 7297 10659
rect 7331 10625 7343 10659
rect 7285 10619 7343 10625
rect 5902 10548 5908 10600
rect 5960 10588 5966 10600
rect 6270 10588 6276 10600
rect 5960 10560 6276 10588
rect 5960 10548 5966 10560
rect 6270 10548 6276 10560
rect 6328 10548 6334 10600
rect 6365 10591 6423 10597
rect 6365 10557 6377 10591
rect 6411 10588 6423 10591
rect 7098 10588 7104 10600
rect 6411 10560 7104 10588
rect 6411 10557 6423 10560
rect 6365 10551 6423 10557
rect 6380 10452 6408 10551
rect 7098 10548 7104 10560
rect 7156 10548 7162 10600
rect 12342 10548 12348 10600
rect 12400 10588 12406 10600
rect 12544 10597 12572 10696
rect 12989 10693 13001 10696
rect 13035 10693 13047 10727
rect 13538 10724 13544 10736
rect 12989 10687 13047 10693
rect 13372 10696 13544 10724
rect 12710 10616 12716 10668
rect 12768 10616 12774 10668
rect 12897 10659 12955 10665
rect 12897 10625 12909 10659
rect 12943 10656 12955 10659
rect 13372 10656 13400 10696
rect 13538 10684 13544 10696
rect 13596 10724 13602 10736
rect 13596 10696 13676 10724
rect 13596 10684 13602 10696
rect 13648 10665 13676 10696
rect 15654 10684 15660 10736
rect 15712 10684 15718 10736
rect 12943 10628 13400 10656
rect 13449 10659 13507 10665
rect 12943 10625 12955 10628
rect 12897 10619 12955 10625
rect 13449 10625 13461 10659
rect 13495 10625 13507 10659
rect 13449 10619 13507 10625
rect 13633 10659 13691 10665
rect 13633 10625 13645 10659
rect 13679 10625 13691 10659
rect 13633 10619 13691 10625
rect 12529 10591 12587 10597
rect 12529 10588 12541 10591
rect 12400 10560 12541 10588
rect 12400 10548 12406 10560
rect 12529 10557 12541 10560
rect 12575 10557 12587 10591
rect 12529 10551 12587 10557
rect 13354 10548 13360 10600
rect 13412 10588 13418 10600
rect 13464 10588 13492 10619
rect 13412 10560 13492 10588
rect 13412 10548 13418 10560
rect 13541 10523 13599 10529
rect 13541 10520 13553 10523
rect 13188 10492 13553 10520
rect 5736 10424 6408 10452
rect 7469 10455 7527 10461
rect 7469 10421 7481 10455
rect 7515 10452 7527 10455
rect 7742 10452 7748 10464
rect 7515 10424 7748 10452
rect 7515 10421 7527 10424
rect 7469 10415 7527 10421
rect 7742 10412 7748 10424
rect 7800 10452 7806 10464
rect 8294 10452 8300 10464
rect 7800 10424 8300 10452
rect 7800 10412 7806 10424
rect 8294 10412 8300 10424
rect 8352 10412 8358 10464
rect 8386 10412 8392 10464
rect 8444 10452 8450 10464
rect 9306 10452 9312 10464
rect 8444 10424 9312 10452
rect 8444 10412 8450 10424
rect 9306 10412 9312 10424
rect 9364 10412 9370 10464
rect 13188 10461 13216 10492
rect 13541 10489 13553 10492
rect 13587 10489 13599 10523
rect 13541 10483 13599 10489
rect 13173 10455 13231 10461
rect 13173 10421 13185 10455
rect 13219 10421 13231 10455
rect 13173 10415 13231 10421
rect 1104 10362 16376 10384
rect 1104 10310 2859 10362
rect 2911 10310 2923 10362
rect 2975 10310 2987 10362
rect 3039 10310 3051 10362
rect 3103 10310 3115 10362
rect 3167 10310 6677 10362
rect 6729 10310 6741 10362
rect 6793 10310 6805 10362
rect 6857 10310 6869 10362
rect 6921 10310 6933 10362
rect 6985 10310 10495 10362
rect 10547 10310 10559 10362
rect 10611 10310 10623 10362
rect 10675 10310 10687 10362
rect 10739 10310 10751 10362
rect 10803 10310 14313 10362
rect 14365 10310 14377 10362
rect 14429 10310 14441 10362
rect 14493 10310 14505 10362
rect 14557 10310 14569 10362
rect 14621 10310 16376 10362
rect 1104 10288 16376 10310
rect 2406 10208 2412 10260
rect 2464 10248 2470 10260
rect 3421 10251 3479 10257
rect 2464 10220 2774 10248
rect 2464 10208 2470 10220
rect 2746 10112 2774 10220
rect 3421 10217 3433 10251
rect 3467 10248 3479 10251
rect 3878 10248 3884 10260
rect 3467 10220 3884 10248
rect 3467 10217 3479 10220
rect 3421 10211 3479 10217
rect 3878 10208 3884 10220
rect 3936 10208 3942 10260
rect 5169 10251 5227 10257
rect 5169 10248 5181 10251
rect 4172 10220 5181 10248
rect 3602 10140 3608 10192
rect 3660 10180 3666 10192
rect 4172 10180 4200 10220
rect 5169 10217 5181 10220
rect 5215 10217 5227 10251
rect 5169 10211 5227 10217
rect 5534 10208 5540 10260
rect 5592 10248 5598 10260
rect 5994 10248 6000 10260
rect 5592 10220 6000 10248
rect 5592 10208 5598 10220
rect 5994 10208 6000 10220
rect 6052 10208 6058 10260
rect 6086 10208 6092 10260
rect 6144 10248 6150 10260
rect 6365 10251 6423 10257
rect 6365 10248 6377 10251
rect 6144 10220 6377 10248
rect 6144 10208 6150 10220
rect 6365 10217 6377 10220
rect 6411 10217 6423 10251
rect 6365 10211 6423 10217
rect 8297 10251 8355 10257
rect 8297 10217 8309 10251
rect 8343 10248 8355 10251
rect 8386 10248 8392 10260
rect 8343 10220 8392 10248
rect 8343 10217 8355 10220
rect 8297 10211 8355 10217
rect 8386 10208 8392 10220
rect 8444 10248 8450 10260
rect 9490 10248 9496 10260
rect 8444 10220 9496 10248
rect 8444 10208 8450 10220
rect 9490 10208 9496 10220
rect 9548 10208 9554 10260
rect 9585 10251 9643 10257
rect 9585 10217 9597 10251
rect 9631 10248 9643 10251
rect 9631 10220 11836 10248
rect 9631 10217 9643 10220
rect 9585 10211 9643 10217
rect 3660 10152 4200 10180
rect 3660 10140 3666 10152
rect 4338 10140 4344 10192
rect 4396 10140 4402 10192
rect 4908 10152 5672 10180
rect 4356 10112 4384 10140
rect 2746 10084 4016 10112
rect 4356 10084 4568 10112
rect 1765 10047 1823 10053
rect 1765 10013 1777 10047
rect 1811 10044 1823 10047
rect 1811 10016 2774 10044
rect 1811 10013 1823 10016
rect 1765 10007 1823 10013
rect 1486 9868 1492 9920
rect 1544 9868 1550 9920
rect 2746 9908 2774 10016
rect 3234 10004 3240 10056
rect 3292 10044 3298 10056
rect 3436 10053 3464 10084
rect 3988 10053 4016 10084
rect 3421 10047 3479 10053
rect 3292 10016 3372 10044
rect 3292 10004 3298 10016
rect 3344 9976 3372 10016
rect 3421 10013 3433 10047
rect 3467 10013 3479 10047
rect 3421 10007 3479 10013
rect 3789 10047 3847 10053
rect 3789 10013 3801 10047
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 3973 10047 4031 10053
rect 3973 10013 3985 10047
rect 4019 10013 4031 10047
rect 3973 10007 4031 10013
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10044 4215 10047
rect 4249 10047 4307 10053
rect 4249 10044 4261 10047
rect 4203 10016 4261 10044
rect 4203 10013 4215 10016
rect 4157 10007 4215 10013
rect 4249 10013 4261 10016
rect 4295 10013 4307 10047
rect 4249 10007 4307 10013
rect 3804 9976 3832 10007
rect 4430 10004 4436 10056
rect 4488 10004 4494 10056
rect 4540 10053 4568 10084
rect 4525 10047 4583 10053
rect 4525 10013 4537 10047
rect 4571 10013 4583 10047
rect 4525 10007 4583 10013
rect 4614 10004 4620 10056
rect 4672 10044 4678 10056
rect 4908 10053 4936 10152
rect 5644 10124 5672 10152
rect 5902 10140 5908 10192
rect 5960 10180 5966 10192
rect 9674 10180 9680 10192
rect 5960 10152 9680 10180
rect 5960 10140 5966 10152
rect 9674 10140 9680 10152
rect 9732 10140 9738 10192
rect 9861 10183 9919 10189
rect 9861 10149 9873 10183
rect 9907 10180 9919 10183
rect 9950 10180 9956 10192
rect 9907 10152 9956 10180
rect 9907 10149 9919 10152
rect 9861 10143 9919 10149
rect 9950 10140 9956 10152
rect 10008 10140 10014 10192
rect 4985 10115 5043 10121
rect 4985 10081 4997 10115
rect 5031 10112 5043 10115
rect 5031 10084 5212 10112
rect 5031 10081 5043 10084
rect 4985 10075 5043 10081
rect 4709 10047 4767 10053
rect 4709 10044 4721 10047
rect 4672 10016 4721 10044
rect 4672 10004 4678 10016
rect 4709 10013 4721 10016
rect 4755 10013 4767 10047
rect 4709 10007 4767 10013
rect 4893 10047 4951 10053
rect 4893 10013 4905 10047
rect 4939 10013 4951 10047
rect 4893 10007 4951 10013
rect 5074 10004 5080 10056
rect 5132 10004 5138 10056
rect 5184 10053 5212 10084
rect 5626 10072 5632 10124
rect 5684 10072 5690 10124
rect 6362 10112 6368 10124
rect 5920 10084 6368 10112
rect 5169 10047 5227 10053
rect 5169 10013 5181 10047
rect 5215 10013 5227 10047
rect 5169 10007 5227 10013
rect 5353 10047 5411 10053
rect 5353 10013 5365 10047
rect 5399 10044 5411 10047
rect 5718 10044 5724 10056
rect 5399 10016 5724 10044
rect 5399 10013 5411 10016
rect 5353 10007 5411 10013
rect 5718 10004 5724 10016
rect 5776 10004 5782 10056
rect 5810 10004 5816 10056
rect 5868 10044 5874 10056
rect 5920 10053 5948 10084
rect 6362 10072 6368 10084
rect 6420 10112 6426 10124
rect 9125 10115 9183 10121
rect 6420 10084 6776 10112
rect 6420 10072 6426 10084
rect 5905 10047 5963 10053
rect 5905 10044 5917 10047
rect 5868 10016 5917 10044
rect 5868 10004 5874 10016
rect 5905 10013 5917 10016
rect 5951 10013 5963 10047
rect 5905 10007 5963 10013
rect 6086 10004 6092 10056
rect 6144 10004 6150 10056
rect 6454 10004 6460 10056
rect 6512 10004 6518 10056
rect 6546 10004 6552 10056
rect 6604 10004 6610 10056
rect 6748 10053 6776 10084
rect 9125 10081 9137 10115
rect 9171 10112 9183 10115
rect 10321 10115 10379 10121
rect 10321 10112 10333 10115
rect 9171 10084 10333 10112
rect 9171 10081 9183 10084
rect 9125 10075 9183 10081
rect 10321 10081 10333 10084
rect 10367 10081 10379 10115
rect 11808 10112 11836 10220
rect 12342 10208 12348 10260
rect 12400 10208 12406 10260
rect 12710 10208 12716 10260
rect 12768 10208 12774 10260
rect 14826 10208 14832 10260
rect 14884 10248 14890 10260
rect 14921 10251 14979 10257
rect 14921 10248 14933 10251
rect 14884 10220 14933 10248
rect 14884 10208 14890 10220
rect 14921 10217 14933 10220
rect 14967 10217 14979 10251
rect 14921 10211 14979 10217
rect 11808 10084 12204 10112
rect 10321 10075 10379 10081
rect 6733 10047 6791 10053
rect 6733 10013 6745 10047
rect 6779 10013 6791 10047
rect 6733 10007 6791 10013
rect 6914 10004 6920 10056
rect 6972 10004 6978 10056
rect 9030 10004 9036 10056
rect 9088 10044 9094 10056
rect 9217 10047 9275 10053
rect 9217 10044 9229 10047
rect 9088 10016 9229 10044
rect 9088 10004 9094 10016
rect 9217 10013 9229 10016
rect 9263 10013 9275 10047
rect 9217 10007 9275 10013
rect 9306 10004 9312 10056
rect 9364 10004 9370 10056
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10013 9459 10047
rect 9401 10007 9459 10013
rect 6472 9976 6500 10004
rect 6641 9979 6699 9985
rect 6641 9976 6653 9979
rect 3344 9948 3832 9976
rect 4356 9948 6224 9976
rect 6472 9948 6653 9976
rect 4154 9908 4160 9920
rect 2746 9880 4160 9908
rect 4154 9868 4160 9880
rect 4212 9868 4218 9920
rect 4356 9917 4384 9948
rect 4341 9911 4399 9917
rect 4341 9877 4353 9911
rect 4387 9877 4399 9911
rect 4341 9871 4399 9877
rect 4709 9911 4767 9917
rect 4709 9877 4721 9911
rect 4755 9908 4767 9911
rect 5902 9908 5908 9920
rect 4755 9880 5908 9908
rect 4755 9877 4767 9880
rect 4709 9871 4767 9877
rect 5902 9868 5908 9880
rect 5960 9868 5966 9920
rect 6196 9908 6224 9948
rect 6641 9945 6653 9948
rect 6687 9945 6699 9979
rect 6641 9939 6699 9945
rect 8110 9936 8116 9988
rect 8168 9936 8174 9988
rect 8329 9979 8387 9985
rect 8329 9945 8341 9979
rect 8375 9976 8387 9979
rect 8570 9976 8576 9988
rect 8375 9948 8576 9976
rect 8375 9945 8387 9948
rect 8329 9939 8387 9945
rect 8570 9936 8576 9948
rect 8628 9936 8634 9988
rect 8202 9908 8208 9920
rect 6196 9880 8208 9908
rect 8202 9868 8208 9880
rect 8260 9868 8266 9920
rect 8481 9911 8539 9917
rect 8481 9877 8493 9911
rect 8527 9908 8539 9911
rect 9416 9908 9444 10007
rect 9490 10004 9496 10056
rect 9548 10044 9554 10056
rect 9677 10047 9735 10053
rect 9677 10044 9689 10047
rect 9548 10016 9689 10044
rect 9548 10004 9554 10016
rect 9677 10013 9689 10016
rect 9723 10013 9735 10047
rect 9677 10007 9735 10013
rect 9950 10004 9956 10056
rect 10008 10044 10014 10056
rect 10137 10047 10195 10053
rect 10137 10044 10149 10047
rect 10008 10016 10149 10044
rect 10008 10004 10014 10016
rect 10137 10013 10149 10016
rect 10183 10044 10195 10047
rect 10229 10047 10287 10053
rect 10229 10044 10241 10047
rect 10183 10016 10241 10044
rect 10183 10013 10195 10016
rect 10137 10007 10195 10013
rect 10229 10013 10241 10016
rect 10275 10013 10287 10047
rect 10229 10007 10287 10013
rect 10413 10047 10471 10053
rect 10413 10013 10425 10047
rect 10459 10013 10471 10047
rect 10413 10007 10471 10013
rect 11885 10047 11943 10053
rect 11885 10013 11897 10047
rect 11931 10044 11943 10047
rect 12066 10044 12072 10056
rect 11931 10016 12072 10044
rect 11931 10013 11943 10016
rect 11885 10007 11943 10013
rect 10318 9976 10324 9988
rect 10060 9948 10324 9976
rect 10060 9917 10088 9948
rect 10318 9936 10324 9948
rect 10376 9976 10382 9988
rect 10428 9976 10456 10007
rect 12066 10004 12072 10016
rect 12124 10004 12130 10056
rect 12176 10053 12204 10084
rect 12161 10047 12219 10053
rect 12161 10013 12173 10047
rect 12207 10044 12219 10047
rect 12437 10047 12495 10053
rect 12437 10044 12449 10047
rect 12207 10016 12449 10044
rect 12207 10013 12219 10016
rect 12161 10007 12219 10013
rect 12437 10013 12449 10016
rect 12483 10013 12495 10047
rect 12713 10047 12771 10053
rect 12713 10044 12725 10047
rect 12437 10007 12495 10013
rect 12544 10016 12725 10044
rect 12544 9976 12572 10016
rect 12713 10013 12725 10016
rect 12759 10013 12771 10047
rect 12713 10007 12771 10013
rect 14826 10004 14832 10056
rect 14884 10044 14890 10056
rect 15105 10047 15163 10053
rect 15105 10044 15117 10047
rect 14884 10016 15117 10044
rect 14884 10004 14890 10016
rect 15105 10013 15117 10016
rect 15151 10013 15163 10047
rect 15105 10007 15163 10013
rect 15381 10047 15439 10053
rect 15381 10013 15393 10047
rect 15427 10044 15439 10047
rect 15427 10016 15608 10044
rect 15427 10013 15439 10016
rect 15381 10007 15439 10013
rect 10376 9948 10456 9976
rect 12176 9948 12572 9976
rect 12621 9979 12679 9985
rect 10376 9936 10382 9948
rect 10045 9911 10103 9917
rect 10045 9908 10057 9911
rect 8527 9880 10057 9908
rect 8527 9877 8539 9880
rect 8481 9871 8539 9877
rect 10045 9877 10057 9880
rect 10091 9877 10103 9911
rect 10045 9871 10103 9877
rect 11514 9868 11520 9920
rect 11572 9908 11578 9920
rect 11977 9911 12035 9917
rect 11977 9908 11989 9911
rect 11572 9880 11989 9908
rect 11572 9868 11578 9880
rect 11977 9877 11989 9880
rect 12023 9908 12035 9911
rect 12176 9908 12204 9948
rect 12621 9945 12633 9979
rect 12667 9945 12679 9979
rect 12621 9939 12679 9945
rect 12023 9880 12204 9908
rect 12023 9877 12035 9880
rect 11977 9871 12035 9877
rect 12250 9868 12256 9920
rect 12308 9908 12314 9920
rect 12636 9908 12664 9939
rect 15580 9920 15608 10016
rect 15654 9936 15660 9988
rect 15712 9936 15718 9988
rect 12308 9880 12664 9908
rect 15289 9911 15347 9917
rect 12308 9868 12314 9880
rect 15289 9877 15301 9911
rect 15335 9908 15347 9911
rect 15378 9908 15384 9920
rect 15335 9880 15384 9908
rect 15335 9877 15347 9880
rect 15289 9871 15347 9877
rect 15378 9868 15384 9880
rect 15436 9868 15442 9920
rect 15562 9868 15568 9920
rect 15620 9868 15626 9920
rect 15933 9911 15991 9917
rect 15933 9877 15945 9911
rect 15979 9908 15991 9911
rect 16022 9908 16028 9920
rect 15979 9880 16028 9908
rect 15979 9877 15991 9880
rect 15933 9871 15991 9877
rect 16022 9868 16028 9880
rect 16080 9868 16086 9920
rect 1104 9818 16376 9840
rect 1104 9766 3519 9818
rect 3571 9766 3583 9818
rect 3635 9766 3647 9818
rect 3699 9766 3711 9818
rect 3763 9766 3775 9818
rect 3827 9766 7337 9818
rect 7389 9766 7401 9818
rect 7453 9766 7465 9818
rect 7517 9766 7529 9818
rect 7581 9766 7593 9818
rect 7645 9766 11155 9818
rect 11207 9766 11219 9818
rect 11271 9766 11283 9818
rect 11335 9766 11347 9818
rect 11399 9766 11411 9818
rect 11463 9766 14973 9818
rect 15025 9766 15037 9818
rect 15089 9766 15101 9818
rect 15153 9766 15165 9818
rect 15217 9766 15229 9818
rect 15281 9766 16376 9818
rect 1104 9744 16376 9766
rect 3145 9707 3203 9713
rect 3145 9673 3157 9707
rect 3191 9704 3203 9707
rect 3234 9704 3240 9716
rect 3191 9676 3240 9704
rect 3191 9673 3203 9676
rect 3145 9667 3203 9673
rect 3234 9664 3240 9676
rect 3292 9664 3298 9716
rect 3418 9664 3424 9716
rect 3476 9704 3482 9716
rect 7006 9704 7012 9716
rect 3476 9676 7012 9704
rect 3476 9664 3482 9676
rect 7006 9664 7012 9676
rect 7064 9664 7070 9716
rect 7653 9707 7711 9713
rect 7300 9676 7512 9704
rect 4157 9639 4215 9645
rect 4157 9636 4169 9639
rect 3068 9608 4169 9636
rect 1670 9528 1676 9580
rect 1728 9568 1734 9580
rect 3068 9577 3096 9608
rect 4157 9605 4169 9608
rect 4203 9605 4215 9639
rect 4338 9636 4344 9648
rect 4157 9599 4215 9605
rect 4264 9608 4344 9636
rect 3053 9571 3111 9577
rect 3053 9568 3065 9571
rect 1728 9540 3065 9568
rect 1728 9528 1734 9540
rect 3053 9537 3065 9540
rect 3099 9537 3111 9571
rect 3053 9531 3111 9537
rect 3237 9571 3295 9577
rect 3237 9537 3249 9571
rect 3283 9537 3295 9571
rect 3237 9531 3295 9537
rect 3252 9500 3280 9531
rect 3326 9528 3332 9580
rect 3384 9568 3390 9580
rect 3513 9571 3571 9577
rect 3513 9568 3525 9571
rect 3384 9540 3525 9568
rect 3384 9528 3390 9540
rect 3513 9537 3525 9540
rect 3559 9537 3571 9571
rect 3513 9531 3571 9537
rect 3697 9571 3755 9577
rect 3697 9537 3709 9571
rect 3743 9568 3755 9571
rect 3973 9571 4031 9577
rect 3973 9568 3985 9571
rect 3743 9540 3985 9568
rect 3743 9537 3755 9540
rect 3697 9531 3755 9537
rect 3973 9537 3985 9540
rect 4019 9537 4031 9571
rect 4264 9568 4292 9608
rect 4338 9596 4344 9608
rect 4396 9596 4402 9648
rect 4522 9596 4528 9648
rect 4580 9636 4586 9648
rect 6914 9636 6920 9648
rect 4580 9608 6920 9636
rect 4580 9596 4586 9608
rect 6914 9596 6920 9608
rect 6972 9596 6978 9648
rect 7300 9636 7328 9676
rect 7116 9608 7328 9636
rect 7484 9636 7512 9676
rect 7653 9673 7665 9707
rect 7699 9673 7711 9707
rect 7653 9667 7711 9673
rect 7558 9636 7564 9648
rect 7484 9608 7564 9636
rect 7116 9577 7144 9608
rect 7558 9596 7564 9608
rect 7616 9596 7622 9648
rect 7668 9636 7696 9667
rect 8202 9664 8208 9716
rect 8260 9704 8266 9716
rect 8260 9676 13308 9704
rect 8260 9664 8266 9676
rect 8110 9636 8116 9648
rect 7668 9608 8116 9636
rect 8110 9596 8116 9608
rect 8168 9636 8174 9648
rect 8297 9639 8355 9645
rect 8297 9636 8309 9639
rect 8168 9608 8309 9636
rect 8168 9596 8174 9608
rect 8297 9605 8309 9608
rect 8343 9605 8355 9639
rect 8297 9599 8355 9605
rect 8386 9596 8392 9648
rect 8444 9596 8450 9648
rect 8481 9639 8539 9645
rect 8481 9605 8493 9639
rect 8527 9636 8539 9639
rect 8570 9636 8576 9648
rect 8527 9608 8576 9636
rect 8527 9605 8539 9608
rect 8481 9599 8539 9605
rect 8570 9596 8576 9608
rect 8628 9596 8634 9648
rect 9030 9596 9036 9648
rect 9088 9596 9094 9648
rect 11149 9639 11207 9645
rect 9263 9605 9321 9611
rect 9263 9602 9275 9605
rect 3973 9531 4031 9537
rect 4080 9540 4292 9568
rect 7101 9571 7159 9577
rect 4080 9500 4108 9540
rect 7101 9537 7113 9571
rect 7147 9537 7159 9571
rect 7101 9531 7159 9537
rect 7285 9571 7343 9577
rect 7285 9537 7297 9571
rect 7331 9537 7343 9571
rect 7285 9531 7343 9537
rect 3252 9472 4108 9500
rect 7190 9460 7196 9512
rect 7248 9500 7254 9512
rect 7300 9500 7328 9531
rect 7374 9528 7380 9580
rect 7432 9528 7438 9580
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9568 7527 9571
rect 7650 9568 7656 9580
rect 7515 9540 7656 9568
rect 7515 9537 7527 9540
rect 7469 9531 7527 9537
rect 7650 9528 7656 9540
rect 7708 9528 7714 9580
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9537 7803 9571
rect 7745 9531 7803 9537
rect 8205 9571 8263 9577
rect 8205 9537 8217 9571
rect 8251 9568 8263 9571
rect 8404 9568 8432 9596
rect 8251 9540 8432 9568
rect 8251 9537 8263 9540
rect 8205 9531 8263 9537
rect 7248 9472 7328 9500
rect 7248 9460 7254 9472
rect 7466 9392 7472 9444
rect 7524 9432 7530 9444
rect 7760 9432 7788 9531
rect 7837 9503 7895 9509
rect 7837 9469 7849 9503
rect 7883 9469 7895 9503
rect 7837 9463 7895 9469
rect 7524 9404 7788 9432
rect 7524 9392 7530 9404
rect 3878 9324 3884 9376
rect 3936 9324 3942 9376
rect 6454 9324 6460 9376
rect 6512 9364 6518 9376
rect 7852 9364 7880 9463
rect 8113 9435 8171 9441
rect 8113 9401 8125 9435
rect 8159 9432 8171 9435
rect 8220 9432 8248 9531
rect 9122 9528 9128 9580
rect 9180 9568 9186 9580
rect 9248 9571 9275 9602
rect 9309 9571 9321 9605
rect 10336 9608 10916 9636
rect 10336 9580 10364 9608
rect 9248 9568 9321 9571
rect 9180 9565 9321 9568
rect 9180 9540 9276 9565
rect 9180 9528 9186 9540
rect 10318 9528 10324 9580
rect 10376 9528 10382 9580
rect 10888 9577 10916 9608
rect 11149 9605 11161 9639
rect 11195 9605 11207 9639
rect 13280 9636 13308 9676
rect 13354 9664 13360 9716
rect 13412 9664 13418 9716
rect 13906 9704 13912 9716
rect 13464 9676 13912 9704
rect 13464 9636 13492 9676
rect 13906 9664 13912 9676
rect 13964 9664 13970 9716
rect 13280 9608 13492 9636
rect 11149 9599 11207 9605
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9537 10471 9571
rect 10413 9531 10471 9537
rect 10873 9571 10931 9577
rect 10873 9537 10885 9571
rect 10919 9537 10931 9571
rect 11164 9568 11192 9599
rect 11701 9571 11759 9577
rect 11701 9568 11713 9571
rect 11164 9540 11713 9568
rect 10873 9531 10931 9537
rect 11701 9537 11713 9540
rect 11747 9537 11759 9571
rect 11701 9531 11759 9537
rect 10428 9500 10456 9531
rect 13170 9528 13176 9580
rect 13228 9568 13234 9580
rect 13541 9571 13599 9577
rect 13541 9568 13553 9571
rect 13228 9540 13553 9568
rect 13228 9528 13234 9540
rect 13541 9537 13553 9540
rect 13587 9537 13599 9571
rect 13541 9531 13599 9537
rect 13630 9528 13636 9580
rect 13688 9568 13694 9580
rect 13725 9571 13783 9577
rect 13725 9568 13737 9571
rect 13688 9540 13737 9568
rect 13688 9528 13694 9540
rect 13725 9537 13737 9540
rect 13771 9537 13783 9571
rect 13725 9531 13783 9537
rect 13998 9528 14004 9580
rect 14056 9568 14062 9580
rect 14642 9568 14648 9580
rect 14056 9540 14648 9568
rect 14056 9528 14062 9540
rect 14642 9528 14648 9540
rect 14700 9568 14706 9580
rect 14829 9571 14887 9577
rect 14829 9568 14841 9571
rect 14700 9540 14841 9568
rect 14700 9528 14706 9540
rect 14829 9537 14841 9540
rect 14875 9537 14887 9571
rect 14829 9531 14887 9537
rect 15378 9528 15384 9580
rect 15436 9568 15442 9580
rect 15473 9571 15531 9577
rect 15473 9568 15485 9571
rect 15436 9540 15485 9568
rect 15436 9528 15442 9540
rect 15473 9537 15485 9540
rect 15519 9537 15531 9571
rect 15473 9531 15531 9537
rect 8496 9472 10456 9500
rect 8496 9441 8524 9472
rect 8159 9404 8248 9432
rect 8481 9435 8539 9441
rect 8159 9401 8171 9404
rect 8113 9395 8171 9401
rect 8481 9401 8493 9435
rect 8527 9401 8539 9435
rect 8481 9395 8539 9401
rect 9401 9435 9459 9441
rect 9401 9401 9413 9435
rect 9447 9432 9459 9435
rect 9950 9432 9956 9444
rect 9447 9404 9956 9432
rect 9447 9401 9459 9404
rect 9401 9395 9459 9401
rect 9950 9392 9956 9404
rect 10008 9392 10014 9444
rect 10428 9432 10456 9472
rect 10502 9460 10508 9512
rect 10560 9500 10566 9512
rect 11149 9503 11207 9509
rect 11149 9500 11161 9503
rect 10560 9472 11161 9500
rect 10560 9460 10566 9472
rect 11149 9469 11161 9472
rect 11195 9469 11207 9503
rect 11514 9500 11520 9512
rect 11149 9463 11207 9469
rect 11440 9472 11520 9500
rect 10965 9435 11023 9441
rect 10965 9432 10977 9435
rect 10428 9404 10977 9432
rect 10965 9401 10977 9404
rect 11011 9401 11023 9435
rect 10965 9395 11023 9401
rect 6512 9336 7880 9364
rect 7929 9367 7987 9373
rect 6512 9324 6518 9336
rect 7929 9333 7941 9367
rect 7975 9364 7987 9367
rect 8018 9364 8024 9376
rect 7975 9336 8024 9364
rect 7975 9333 7987 9336
rect 7929 9327 7987 9333
rect 8018 9324 8024 9336
rect 8076 9324 8082 9376
rect 9217 9367 9275 9373
rect 9217 9333 9229 9367
rect 9263 9364 9275 9367
rect 9306 9364 9312 9376
rect 9263 9336 9312 9364
rect 9263 9333 9275 9336
rect 9217 9327 9275 9333
rect 9306 9324 9312 9336
rect 9364 9324 9370 9376
rect 10318 9324 10324 9376
rect 10376 9364 10382 9376
rect 10413 9367 10471 9373
rect 10413 9364 10425 9367
rect 10376 9336 10425 9364
rect 10376 9324 10382 9336
rect 10413 9333 10425 9336
rect 10459 9333 10471 9367
rect 10413 9327 10471 9333
rect 10781 9367 10839 9373
rect 10781 9333 10793 9367
rect 10827 9364 10839 9367
rect 11440 9364 11468 9472
rect 11514 9460 11520 9472
rect 11572 9460 11578 9512
rect 12989 9503 13047 9509
rect 12989 9469 13001 9503
rect 13035 9500 13047 9503
rect 13648 9500 13676 9528
rect 13035 9472 13676 9500
rect 14553 9503 14611 9509
rect 13035 9469 13047 9472
rect 12989 9463 13047 9469
rect 14553 9469 14565 9503
rect 14599 9500 14611 9503
rect 14734 9500 14740 9512
rect 14599 9472 14740 9500
rect 14599 9469 14611 9472
rect 14553 9463 14611 9469
rect 14734 9460 14740 9472
rect 14792 9460 14798 9512
rect 15197 9503 15255 9509
rect 15197 9469 15209 9503
rect 15243 9500 15255 9503
rect 15562 9500 15568 9512
rect 15243 9472 15568 9500
rect 15243 9469 15255 9472
rect 15197 9463 15255 9469
rect 15562 9460 15568 9472
rect 15620 9460 15626 9512
rect 15654 9460 15660 9512
rect 15712 9500 15718 9512
rect 15841 9503 15899 9509
rect 15841 9500 15853 9503
rect 15712 9472 15853 9500
rect 15712 9460 15718 9472
rect 15841 9469 15853 9472
rect 15887 9469 15899 9503
rect 15841 9463 15899 9469
rect 10827 9336 11468 9364
rect 10827 9333 10839 9336
rect 10781 9327 10839 9333
rect 11882 9324 11888 9376
rect 11940 9324 11946 9376
rect 1104 9274 16376 9296
rect 1104 9222 2859 9274
rect 2911 9222 2923 9274
rect 2975 9222 2987 9274
rect 3039 9222 3051 9274
rect 3103 9222 3115 9274
rect 3167 9222 6677 9274
rect 6729 9222 6741 9274
rect 6793 9222 6805 9274
rect 6857 9222 6869 9274
rect 6921 9222 6933 9274
rect 6985 9222 10495 9274
rect 10547 9222 10559 9274
rect 10611 9222 10623 9274
rect 10675 9222 10687 9274
rect 10739 9222 10751 9274
rect 10803 9222 14313 9274
rect 14365 9222 14377 9274
rect 14429 9222 14441 9274
rect 14493 9222 14505 9274
rect 14557 9222 14569 9274
rect 14621 9222 16376 9274
rect 1104 9200 16376 9222
rect 4338 9120 4344 9172
rect 4396 9160 4402 9172
rect 4709 9163 4767 9169
rect 4709 9160 4721 9163
rect 4396 9132 4721 9160
rect 4396 9120 4402 9132
rect 4709 9129 4721 9132
rect 4755 9129 4767 9163
rect 4709 9123 4767 9129
rect 5445 9163 5503 9169
rect 5445 9129 5457 9163
rect 5491 9129 5503 9163
rect 5445 9123 5503 9129
rect 7009 9163 7067 9169
rect 7009 9129 7021 9163
rect 7055 9160 7067 9163
rect 9766 9160 9772 9172
rect 7055 9132 9772 9160
rect 7055 9129 7067 9132
rect 7009 9123 7067 9129
rect 5261 9095 5319 9101
rect 5261 9061 5273 9095
rect 5307 9061 5319 9095
rect 5460 9092 5488 9123
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 11882 9120 11888 9172
rect 11940 9120 11946 9172
rect 12069 9163 12127 9169
rect 12069 9129 12081 9163
rect 12115 9160 12127 9163
rect 12250 9160 12256 9172
rect 12115 9132 12256 9160
rect 12115 9129 12127 9132
rect 12069 9123 12127 9129
rect 12250 9120 12256 9132
rect 12308 9160 12314 9172
rect 12345 9163 12403 9169
rect 12345 9160 12357 9163
rect 12308 9132 12357 9160
rect 12308 9120 12314 9132
rect 12345 9129 12357 9132
rect 12391 9129 12403 9163
rect 12345 9123 12403 9129
rect 13170 9120 13176 9172
rect 13228 9120 13234 9172
rect 14734 9120 14740 9172
rect 14792 9120 14798 9172
rect 14826 9120 14832 9172
rect 14884 9120 14890 9172
rect 5902 9092 5908 9104
rect 5460 9064 5908 9092
rect 5261 9055 5319 9061
rect 5077 9027 5135 9033
rect 5077 8993 5089 9027
rect 5123 9024 5135 9027
rect 5276 9024 5304 9055
rect 5902 9052 5908 9064
rect 5960 9092 5966 9104
rect 6546 9092 6552 9104
rect 5960 9064 6552 9092
rect 5960 9052 5966 9064
rect 5123 8996 5304 9024
rect 5123 8993 5135 8996
rect 5077 8987 5135 8993
rect 6178 8984 6184 9036
rect 6236 8984 6242 9036
rect 4985 8959 5043 8965
rect 4985 8925 4997 8959
rect 5031 8956 5043 8959
rect 5534 8956 5540 8968
rect 5031 8928 5540 8956
rect 5031 8925 5043 8928
rect 4985 8919 5043 8925
rect 5534 8916 5540 8928
rect 5592 8916 5598 8968
rect 5905 8959 5963 8965
rect 5905 8956 5917 8959
rect 5736 8928 5917 8956
rect 5736 8900 5764 8928
rect 5905 8925 5917 8928
rect 5951 8925 5963 8959
rect 5905 8919 5963 8925
rect 6089 8959 6147 8965
rect 6089 8925 6101 8959
rect 6135 8956 6147 8959
rect 6196 8956 6224 8984
rect 6288 8965 6316 9064
rect 6546 9052 6552 9064
rect 6604 9052 6610 9104
rect 7466 9052 7472 9104
rect 7524 9052 7530 9104
rect 8036 9064 8248 9092
rect 7650 9024 7656 9036
rect 7392 8996 7656 9024
rect 6135 8928 6224 8956
rect 6273 8959 6331 8965
rect 6135 8925 6147 8928
rect 6089 8919 6147 8925
rect 6273 8925 6285 8959
rect 6319 8925 6331 8959
rect 6273 8919 6331 8925
rect 6546 8916 6552 8968
rect 6604 8916 6610 8968
rect 6730 8916 6736 8968
rect 6788 8916 6794 8968
rect 7392 8965 7420 8996
rect 7650 8984 7656 8996
rect 7708 9024 7714 9036
rect 8036 9032 8064 9064
rect 7944 9024 8064 9032
rect 7708 9004 8064 9024
rect 7708 8996 7972 9004
rect 7708 8984 7714 8996
rect 8110 8984 8116 9036
rect 8168 8984 8174 9036
rect 8220 9033 8248 9064
rect 8386 9052 8392 9104
rect 8444 9092 8450 9104
rect 9122 9092 9128 9104
rect 8444 9064 9128 9092
rect 8444 9052 8450 9064
rect 9122 9052 9128 9064
rect 9180 9052 9186 9104
rect 11609 9095 11667 9101
rect 11609 9061 11621 9095
rect 11655 9061 11667 9095
rect 11609 9055 11667 9061
rect 8205 9027 8263 9033
rect 8205 8993 8217 9027
rect 8251 8993 8263 9027
rect 9033 9027 9091 9033
rect 9033 9024 9045 9027
rect 8205 8987 8263 8993
rect 8404 8996 9045 9024
rect 8404 8968 8432 8996
rect 9033 8993 9045 8996
rect 9079 8993 9091 9027
rect 9033 8987 9091 8993
rect 7377 8959 7435 8965
rect 7377 8925 7389 8959
rect 7423 8925 7435 8959
rect 7377 8919 7435 8925
rect 7558 8916 7564 8968
rect 7616 8956 7622 8968
rect 8021 8959 8079 8965
rect 7616 8928 7880 8956
rect 7616 8916 7622 8928
rect 934 8848 940 8900
rect 992 8888 998 8900
rect 1397 8891 1455 8897
rect 1397 8888 1409 8891
rect 992 8860 1409 8888
rect 992 8848 998 8860
rect 1397 8857 1409 8860
rect 1443 8857 1455 8891
rect 1397 8851 1455 8857
rect 1762 8848 1768 8900
rect 1820 8848 1826 8900
rect 5629 8891 5687 8897
rect 5629 8857 5641 8891
rect 5675 8888 5687 8891
rect 5718 8888 5724 8900
rect 5675 8860 5724 8888
rect 5675 8857 5687 8860
rect 5629 8851 5687 8857
rect 5718 8848 5724 8860
rect 5776 8848 5782 8900
rect 5994 8848 6000 8900
rect 6052 8888 6058 8900
rect 6181 8891 6239 8897
rect 6181 8888 6193 8891
rect 6052 8860 6193 8888
rect 6052 8848 6058 8860
rect 6181 8857 6193 8860
rect 6227 8857 6239 8891
rect 6564 8888 6592 8916
rect 6181 8851 6239 8857
rect 6288 8860 6592 8888
rect 7101 8891 7159 8897
rect 5429 8823 5487 8829
rect 5429 8789 5441 8823
rect 5475 8820 5487 8823
rect 6288 8820 6316 8860
rect 7101 8857 7113 8891
rect 7147 8857 7159 8891
rect 7101 8851 7159 8857
rect 5475 8792 6316 8820
rect 6457 8823 6515 8829
rect 5475 8789 5487 8792
rect 5429 8783 5487 8789
rect 6457 8789 6469 8823
rect 6503 8820 6515 8823
rect 7116 8820 7144 8851
rect 7852 8832 7880 8928
rect 8021 8925 8033 8959
rect 8067 8956 8079 8959
rect 8297 8959 8355 8965
rect 8067 8928 8248 8956
rect 8067 8925 8079 8928
rect 8021 8919 8079 8925
rect 6503 8792 7144 8820
rect 6503 8789 6515 8792
rect 6457 8783 6515 8789
rect 7834 8780 7840 8832
rect 7892 8780 7898 8832
rect 8220 8820 8248 8928
rect 8297 8925 8309 8959
rect 8343 8956 8355 8959
rect 8386 8956 8392 8968
rect 8343 8928 8392 8956
rect 8343 8925 8355 8928
rect 8297 8919 8355 8925
rect 8386 8916 8392 8928
rect 8444 8916 8450 8968
rect 8570 8916 8576 8968
rect 8628 8916 8634 8968
rect 9140 8965 9168 9052
rect 9493 9027 9551 9033
rect 9493 8993 9505 9027
rect 9539 9024 9551 9027
rect 11624 9024 11652 9055
rect 11900 9024 11928 9120
rect 12158 9052 12164 9104
rect 12216 9092 12222 9104
rect 12216 9064 12848 9092
rect 12216 9052 12222 9064
rect 12820 9033 12848 9064
rect 12253 9027 12311 9033
rect 12253 9024 12265 9027
rect 9539 8996 11468 9024
rect 11624 8996 11836 9024
rect 11900 8996 12265 9024
rect 9539 8993 9551 8996
rect 9493 8987 9551 8993
rect 11440 8965 11468 8996
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8925 9183 8959
rect 9125 8919 9183 8925
rect 11425 8959 11483 8965
rect 11425 8925 11437 8959
rect 11471 8956 11483 8959
rect 11514 8956 11520 8968
rect 11471 8928 11520 8956
rect 11471 8925 11483 8928
rect 11425 8919 11483 8925
rect 11514 8916 11520 8928
rect 11572 8916 11578 8968
rect 11609 8959 11667 8965
rect 11609 8925 11621 8959
rect 11655 8956 11667 8959
rect 11808 8956 11836 8996
rect 12253 8993 12265 8996
rect 12299 8993 12311 9027
rect 12253 8987 12311 8993
rect 12805 9027 12863 9033
rect 12805 8993 12817 9027
rect 12851 8993 12863 9027
rect 12805 8987 12863 8993
rect 11977 8959 12035 8965
rect 11977 8956 11989 8959
rect 11655 8928 11744 8956
rect 11808 8928 11989 8956
rect 11655 8925 11667 8928
rect 11609 8919 11667 8925
rect 8294 8820 8300 8832
rect 8220 8792 8300 8820
rect 8294 8780 8300 8792
rect 8352 8780 8358 8832
rect 8481 8823 8539 8829
rect 8481 8789 8493 8823
rect 8527 8820 8539 8823
rect 8588 8820 8616 8916
rect 11716 8832 11744 8928
rect 11977 8925 11989 8928
rect 12023 8925 12035 8959
rect 12268 8956 12296 8987
rect 12345 8959 12403 8965
rect 12345 8956 12357 8959
rect 12268 8928 12357 8956
rect 11977 8919 12035 8925
rect 12345 8925 12357 8928
rect 12391 8925 12403 8959
rect 12345 8919 12403 8925
rect 12437 8959 12495 8965
rect 12437 8925 12449 8959
rect 12483 8925 12495 8959
rect 12437 8919 12495 8925
rect 12989 8959 13047 8965
rect 12989 8925 13001 8959
rect 13035 8925 13047 8959
rect 12989 8919 13047 8925
rect 11992 8888 12020 8919
rect 12158 8888 12164 8900
rect 11992 8860 12164 8888
rect 12158 8848 12164 8860
rect 12216 8888 12222 8900
rect 12452 8888 12480 8919
rect 13004 8888 13032 8919
rect 14642 8916 14648 8968
rect 14700 8916 14706 8968
rect 14752 8956 14780 9120
rect 14829 8959 14887 8965
rect 14829 8956 14841 8959
rect 14752 8928 14841 8956
rect 14829 8925 14841 8928
rect 14875 8925 14887 8959
rect 14829 8919 14887 8925
rect 12216 8860 12480 8888
rect 12728 8860 13032 8888
rect 12216 8848 12222 8860
rect 8527 8792 8616 8820
rect 8527 8789 8539 8792
rect 8481 8783 8539 8789
rect 11698 8780 11704 8832
rect 11756 8780 11762 8832
rect 12728 8829 12756 8860
rect 12713 8823 12771 8829
rect 12713 8789 12725 8823
rect 12759 8789 12771 8823
rect 12713 8783 12771 8789
rect 1104 8730 16376 8752
rect 1104 8678 3519 8730
rect 3571 8678 3583 8730
rect 3635 8678 3647 8730
rect 3699 8678 3711 8730
rect 3763 8678 3775 8730
rect 3827 8678 7337 8730
rect 7389 8678 7401 8730
rect 7453 8678 7465 8730
rect 7517 8678 7529 8730
rect 7581 8678 7593 8730
rect 7645 8678 11155 8730
rect 11207 8678 11219 8730
rect 11271 8678 11283 8730
rect 11335 8678 11347 8730
rect 11399 8678 11411 8730
rect 11463 8678 14973 8730
rect 15025 8678 15037 8730
rect 15089 8678 15101 8730
rect 15153 8678 15165 8730
rect 15217 8678 15229 8730
rect 15281 8678 16376 8730
rect 1104 8656 16376 8678
rect 3510 8576 3516 8628
rect 3568 8616 3574 8628
rect 3878 8616 3884 8628
rect 3568 8588 3884 8616
rect 3568 8576 3574 8588
rect 3878 8576 3884 8588
rect 3936 8576 3942 8628
rect 5445 8619 5503 8625
rect 5445 8585 5457 8619
rect 5491 8616 5503 8619
rect 5534 8616 5540 8628
rect 5491 8588 5540 8616
rect 5491 8585 5503 8588
rect 5445 8579 5503 8585
rect 5534 8576 5540 8588
rect 5592 8576 5598 8628
rect 5813 8619 5871 8625
rect 5813 8616 5825 8619
rect 5644 8588 5825 8616
rect 5644 8557 5672 8588
rect 5813 8585 5825 8588
rect 5859 8616 5871 8619
rect 6730 8616 6736 8628
rect 5859 8588 6736 8616
rect 5859 8585 5871 8588
rect 5813 8579 5871 8585
rect 6730 8576 6736 8588
rect 6788 8576 6794 8628
rect 7742 8576 7748 8628
rect 7800 8576 7806 8628
rect 8018 8576 8024 8628
rect 8076 8616 8082 8628
rect 8389 8619 8447 8625
rect 8389 8616 8401 8619
rect 8076 8588 8401 8616
rect 8076 8576 8082 8588
rect 8389 8585 8401 8588
rect 8435 8616 8447 8619
rect 9030 8616 9036 8628
rect 8435 8588 9036 8616
rect 8435 8585 8447 8588
rect 8389 8579 8447 8585
rect 9030 8576 9036 8588
rect 9088 8576 9094 8628
rect 9953 8619 10011 8625
rect 9953 8585 9965 8619
rect 9999 8616 10011 8619
rect 10410 8616 10416 8628
rect 9999 8588 10416 8616
rect 9999 8585 10011 8588
rect 9953 8579 10011 8585
rect 10410 8576 10416 8588
rect 10468 8576 10474 8628
rect 11514 8576 11520 8628
rect 11572 8576 11578 8628
rect 12158 8576 12164 8628
rect 12216 8576 12222 8628
rect 15378 8576 15384 8628
rect 15436 8576 15442 8628
rect 3605 8551 3663 8557
rect 3605 8517 3617 8551
rect 3651 8548 3663 8551
rect 5629 8551 5687 8557
rect 3651 8520 4108 8548
rect 3651 8517 3663 8520
rect 3605 8511 3663 8517
rect 4080 8492 4108 8520
rect 5629 8517 5641 8551
rect 5675 8517 5687 8551
rect 5629 8511 5687 8517
rect 6089 8551 6147 8557
rect 6089 8517 6101 8551
rect 6135 8548 6147 8551
rect 6546 8548 6552 8560
rect 6135 8520 6552 8548
rect 6135 8517 6147 8520
rect 6089 8511 6147 8517
rect 2130 8440 2136 8492
rect 2188 8440 2194 8492
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8480 2375 8483
rect 2501 8483 2559 8489
rect 2501 8480 2513 8483
rect 2363 8452 2513 8480
rect 2363 8449 2375 8452
rect 2317 8443 2375 8449
rect 2501 8449 2513 8452
rect 2547 8449 2559 8483
rect 2501 8443 2559 8449
rect 2590 8440 2596 8492
rect 2648 8480 2654 8492
rect 3329 8483 3387 8489
rect 3329 8480 3341 8483
rect 2648 8452 3341 8480
rect 2648 8440 2654 8452
rect 3329 8449 3341 8452
rect 3375 8449 3387 8483
rect 3329 8443 3387 8449
rect 3418 8440 3424 8492
rect 3476 8440 3482 8492
rect 3697 8483 3755 8489
rect 3697 8449 3709 8483
rect 3743 8449 3755 8483
rect 3697 8443 3755 8449
rect 1857 8415 1915 8421
rect 1857 8381 1869 8415
rect 1903 8412 1915 8415
rect 1946 8412 1952 8424
rect 1903 8384 1952 8412
rect 1903 8381 1915 8384
rect 1857 8375 1915 8381
rect 1946 8372 1952 8384
rect 2004 8372 2010 8424
rect 2038 8372 2044 8424
rect 2096 8412 2102 8424
rect 3712 8412 3740 8443
rect 3878 8440 3884 8492
rect 3936 8440 3942 8492
rect 4062 8440 4068 8492
rect 4120 8440 4126 8492
rect 5353 8483 5411 8489
rect 5353 8449 5365 8483
rect 5399 8449 5411 8483
rect 5353 8443 5411 8449
rect 5368 8412 5396 8443
rect 5534 8440 5540 8492
rect 5592 8480 5598 8492
rect 5718 8480 5724 8492
rect 5592 8452 5724 8480
rect 5592 8440 5598 8452
rect 5718 8440 5724 8452
rect 5776 8440 5782 8492
rect 5902 8440 5908 8492
rect 5960 8440 5966 8492
rect 5994 8440 6000 8492
rect 6052 8440 6058 8492
rect 6104 8412 6132 8511
rect 6546 8508 6552 8520
rect 6604 8508 6610 8560
rect 8202 8548 8208 8560
rect 7300 8520 8208 8548
rect 6178 8440 6184 8492
rect 6236 8480 6242 8492
rect 7300 8480 7328 8520
rect 8202 8508 8208 8520
rect 8260 8508 8266 8560
rect 9217 8551 9275 8557
rect 9217 8517 9229 8551
rect 9263 8548 9275 8551
rect 9306 8548 9312 8560
rect 9263 8520 9312 8548
rect 9263 8517 9275 8520
rect 9217 8511 9275 8517
rect 9306 8508 9312 8520
rect 9364 8508 9370 8560
rect 9447 8517 9505 8523
rect 9447 8514 9459 8517
rect 6236 8452 7328 8480
rect 6236 8440 6242 8452
rect 7466 8440 7472 8492
rect 7524 8480 7530 8492
rect 7561 8483 7619 8489
rect 7561 8480 7573 8483
rect 7524 8452 7573 8480
rect 7524 8440 7530 8452
rect 7561 8449 7573 8452
rect 7607 8449 7619 8483
rect 7561 8443 7619 8449
rect 7929 8483 7987 8489
rect 7929 8449 7941 8483
rect 7975 8480 7987 8483
rect 8297 8483 8355 8489
rect 8297 8480 8309 8483
rect 7975 8452 8309 8480
rect 7975 8449 7987 8452
rect 7929 8443 7987 8449
rect 8297 8449 8309 8452
rect 8343 8449 8355 8483
rect 9432 8483 9459 8514
rect 9493 8483 9505 8517
rect 10060 8520 10456 8548
rect 10060 8492 10088 8520
rect 9432 8480 9505 8483
rect 8297 8443 8355 8449
rect 8956 8477 9505 8480
rect 8956 8452 9460 8477
rect 2096 8384 4844 8412
rect 5368 8384 6132 8412
rect 2096 8372 2102 8384
rect 2774 8304 2780 8356
rect 2832 8304 2838 8356
rect 3605 8347 3663 8353
rect 3605 8313 3617 8347
rect 3651 8344 3663 8347
rect 4430 8344 4436 8356
rect 3651 8316 4436 8344
rect 3651 8313 3663 8316
rect 3605 8307 3663 8313
rect 4430 8304 4436 8316
rect 4488 8304 4494 8356
rect 1949 8279 2007 8285
rect 1949 8245 1961 8279
rect 1995 8276 2007 8279
rect 2406 8276 2412 8288
rect 1995 8248 2412 8276
rect 1995 8245 2007 8248
rect 1949 8239 2007 8245
rect 2406 8236 2412 8248
rect 2464 8236 2470 8288
rect 3789 8279 3847 8285
rect 3789 8245 3801 8279
rect 3835 8276 3847 8279
rect 4246 8276 4252 8288
rect 3835 8248 4252 8276
rect 3835 8245 3847 8248
rect 3789 8239 3847 8245
rect 4246 8236 4252 8248
rect 4304 8236 4310 8288
rect 4816 8276 4844 8384
rect 7006 8372 7012 8424
rect 7064 8412 7070 8424
rect 7282 8412 7288 8424
rect 7064 8384 7288 8412
rect 7064 8372 7070 8384
rect 7282 8372 7288 8384
rect 7340 8412 7346 8424
rect 7944 8412 7972 8443
rect 8956 8424 8984 8452
rect 10042 8440 10048 8492
rect 10100 8440 10106 8492
rect 10428 8489 10456 8520
rect 11532 8489 11560 8576
rect 12176 8548 12204 8576
rect 12253 8551 12311 8557
rect 12253 8548 12265 8551
rect 12176 8520 12265 8548
rect 12253 8517 12265 8520
rect 12299 8517 12311 8551
rect 15013 8551 15071 8557
rect 15013 8548 15025 8551
rect 12253 8511 12311 8517
rect 14752 8520 15025 8548
rect 14752 8492 14780 8520
rect 15013 8517 15025 8520
rect 15059 8517 15071 8551
rect 15013 8511 15071 8517
rect 10137 8483 10195 8489
rect 10137 8449 10149 8483
rect 10183 8449 10195 8483
rect 10137 8443 10195 8449
rect 10413 8483 10471 8489
rect 10413 8449 10425 8483
rect 10459 8449 10471 8483
rect 10413 8443 10471 8449
rect 11517 8483 11575 8489
rect 11517 8449 11529 8483
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 7340 8384 7972 8412
rect 7340 8372 7346 8384
rect 8938 8372 8944 8424
rect 8996 8372 9002 8424
rect 9214 8372 9220 8424
rect 9272 8372 9278 8424
rect 9674 8372 9680 8424
rect 9732 8372 9738 8424
rect 10152 8412 10180 8443
rect 11698 8440 11704 8492
rect 11756 8440 11762 8492
rect 11885 8483 11943 8489
rect 11885 8449 11897 8483
rect 11931 8480 11943 8483
rect 12069 8483 12127 8489
rect 12069 8480 12081 8483
rect 11931 8452 12081 8480
rect 11931 8449 11943 8452
rect 11885 8443 11943 8449
rect 12069 8449 12081 8452
rect 12115 8449 12127 8483
rect 12069 8443 12127 8449
rect 14734 8440 14740 8492
rect 14792 8440 14798 8492
rect 14918 8440 14924 8492
rect 14976 8440 14982 8492
rect 15197 8483 15255 8489
rect 15197 8449 15209 8483
rect 15243 8449 15255 8483
rect 15197 8443 15255 8449
rect 10321 8415 10379 8421
rect 10321 8412 10333 8415
rect 10152 8384 10333 8412
rect 5626 8304 5632 8356
rect 5684 8304 5690 8356
rect 7190 8304 7196 8356
rect 7248 8344 7254 8356
rect 8113 8347 8171 8353
rect 8113 8344 8125 8347
rect 7248 8316 8125 8344
rect 7248 8304 7254 8316
rect 8113 8313 8125 8316
rect 8159 8344 8171 8347
rect 9232 8344 9260 8372
rect 9585 8347 9643 8353
rect 8159 8316 9444 8344
rect 8159 8313 8171 8316
rect 8113 8307 8171 8313
rect 7006 8276 7012 8288
rect 4816 8248 7012 8276
rect 7006 8236 7012 8248
rect 7064 8236 7070 8288
rect 9416 8285 9444 8316
rect 9585 8313 9597 8347
rect 9631 8344 9643 8347
rect 10152 8344 10180 8384
rect 10321 8381 10333 8384
rect 10367 8381 10379 8415
rect 10321 8375 10379 8381
rect 9631 8316 10180 8344
rect 10781 8347 10839 8353
rect 9631 8313 9643 8316
rect 9585 8307 9643 8313
rect 10781 8313 10793 8347
rect 10827 8344 10839 8347
rect 11716 8344 11744 8440
rect 14826 8372 14832 8424
rect 14884 8412 14890 8424
rect 15212 8412 15240 8443
rect 14884 8384 15240 8412
rect 14884 8372 14890 8384
rect 10827 8316 11744 8344
rect 10827 8313 10839 8316
rect 10781 8307 10839 8313
rect 9401 8279 9459 8285
rect 9401 8245 9413 8279
rect 9447 8245 9459 8279
rect 9401 8239 9459 8245
rect 12434 8236 12440 8288
rect 12492 8236 12498 8288
rect 1104 8186 16376 8208
rect 1104 8134 2859 8186
rect 2911 8134 2923 8186
rect 2975 8134 2987 8186
rect 3039 8134 3051 8186
rect 3103 8134 3115 8186
rect 3167 8134 6677 8186
rect 6729 8134 6741 8186
rect 6793 8134 6805 8186
rect 6857 8134 6869 8186
rect 6921 8134 6933 8186
rect 6985 8134 10495 8186
rect 10547 8134 10559 8186
rect 10611 8134 10623 8186
rect 10675 8134 10687 8186
rect 10739 8134 10751 8186
rect 10803 8134 14313 8186
rect 14365 8134 14377 8186
rect 14429 8134 14441 8186
rect 14493 8134 14505 8186
rect 14557 8134 14569 8186
rect 14621 8134 16376 8186
rect 1104 8112 16376 8134
rect 1673 8075 1731 8081
rect 1673 8041 1685 8075
rect 1719 8072 1731 8075
rect 1762 8072 1768 8084
rect 1719 8044 1768 8072
rect 1719 8041 1731 8044
rect 1673 8035 1731 8041
rect 1762 8032 1768 8044
rect 1820 8032 1826 8084
rect 1946 8072 1952 8084
rect 1872 8044 1952 8072
rect 1872 7936 1900 8044
rect 1946 8032 1952 8044
rect 2004 8072 2010 8084
rect 2501 8075 2559 8081
rect 2004 8044 2176 8072
rect 2004 8032 2010 8044
rect 2038 7964 2044 8016
rect 2096 7964 2102 8016
rect 1780 7908 1900 7936
rect 1780 7877 1808 7908
rect 1765 7871 1823 7877
rect 1765 7837 1777 7871
rect 1811 7837 1823 7871
rect 1765 7831 1823 7837
rect 1857 7871 1915 7877
rect 1857 7837 1869 7871
rect 1903 7868 1915 7871
rect 2056 7868 2084 7964
rect 2148 7936 2176 8044
rect 2501 8041 2513 8075
rect 2547 8072 2559 8075
rect 2590 8072 2596 8084
rect 2547 8044 2596 8072
rect 2547 8041 2559 8044
rect 2501 8035 2559 8041
rect 2590 8032 2596 8044
rect 2648 8032 2654 8084
rect 2746 8044 4568 8072
rect 2222 7964 2228 8016
rect 2280 8004 2286 8016
rect 2746 8004 2774 8044
rect 2280 7976 2774 8004
rect 4540 8004 4568 8044
rect 4614 8032 4620 8084
rect 4672 8072 4678 8084
rect 5350 8072 5356 8084
rect 4672 8044 5356 8072
rect 4672 8032 4678 8044
rect 5350 8032 5356 8044
rect 5408 8032 5414 8084
rect 7834 8032 7840 8084
rect 7892 8072 7898 8084
rect 8110 8072 8116 8084
rect 7892 8044 8116 8072
rect 7892 8032 7898 8044
rect 8110 8032 8116 8044
rect 8168 8032 8174 8084
rect 8386 8032 8392 8084
rect 8444 8032 8450 8084
rect 8573 8075 8631 8081
rect 8573 8041 8585 8075
rect 8619 8072 8631 8075
rect 8754 8072 8760 8084
rect 8619 8044 8760 8072
rect 8619 8041 8631 8044
rect 8573 8035 8631 8041
rect 8754 8032 8760 8044
rect 8812 8032 8818 8084
rect 12250 8032 12256 8084
rect 12308 8072 12314 8084
rect 12345 8075 12403 8081
rect 12345 8072 12357 8075
rect 12308 8044 12357 8072
rect 12308 8032 12314 8044
rect 12345 8041 12357 8044
rect 12391 8041 12403 8075
rect 12345 8035 12403 8041
rect 14737 8075 14795 8081
rect 14737 8041 14749 8075
rect 14783 8072 14795 8075
rect 14918 8072 14924 8084
rect 14783 8044 14924 8072
rect 14783 8041 14795 8044
rect 14737 8035 14795 8041
rect 5077 8007 5135 8013
rect 5077 8004 5089 8007
rect 4540 7976 5089 8004
rect 2280 7964 2286 7976
rect 5077 7973 5089 7976
rect 5123 8004 5135 8007
rect 5534 8004 5540 8016
rect 5123 7976 5540 8004
rect 5123 7973 5135 7976
rect 5077 7967 5135 7973
rect 5534 7964 5540 7976
rect 5592 7964 5598 8016
rect 6917 8007 6975 8013
rect 6917 7973 6929 8007
rect 6963 8004 6975 8007
rect 8938 8004 8944 8016
rect 6963 7976 8944 8004
rect 6963 7973 6975 7976
rect 6917 7967 6975 7973
rect 8938 7964 8944 7976
rect 8996 8004 9002 8016
rect 9582 8004 9588 8016
rect 8996 7976 9588 8004
rect 8996 7964 9002 7976
rect 9582 7964 9588 7976
rect 9640 7964 9646 8016
rect 12360 8004 12388 8035
rect 14918 8032 14924 8044
rect 14976 8032 14982 8084
rect 13725 8007 13783 8013
rect 12360 7976 12756 8004
rect 2148 7908 2360 7936
rect 1903 7840 2084 7868
rect 1903 7837 1915 7840
rect 1857 7831 1915 7837
rect 1762 7692 1768 7744
rect 1820 7732 1826 7744
rect 1872 7732 1900 7831
rect 2222 7828 2228 7880
rect 2280 7828 2286 7880
rect 2332 7877 2360 7908
rect 2406 7896 2412 7948
rect 2464 7936 2470 7948
rect 3145 7939 3203 7945
rect 3145 7936 3157 7939
rect 2464 7908 3157 7936
rect 2464 7896 2470 7908
rect 3145 7905 3157 7908
rect 3191 7905 3203 7939
rect 3145 7899 3203 7905
rect 3418 7896 3424 7948
rect 3476 7936 3482 7948
rect 3602 7936 3608 7948
rect 3476 7908 3608 7936
rect 3476 7896 3482 7908
rect 3602 7896 3608 7908
rect 3660 7896 3666 7948
rect 4614 7936 4620 7948
rect 4264 7908 4620 7936
rect 2317 7871 2375 7877
rect 2317 7837 2329 7871
rect 2363 7868 2375 7871
rect 2590 7868 2596 7880
rect 2363 7840 2596 7868
rect 2363 7837 2375 7840
rect 2317 7831 2375 7837
rect 2590 7828 2596 7840
rect 2648 7868 2654 7880
rect 2685 7871 2743 7877
rect 2685 7868 2697 7871
rect 2648 7840 2697 7868
rect 2648 7828 2654 7840
rect 2685 7837 2697 7840
rect 2731 7837 2743 7871
rect 2685 7831 2743 7837
rect 3237 7871 3295 7877
rect 3237 7837 3249 7871
rect 3283 7837 3295 7871
rect 3237 7831 3295 7837
rect 2038 7809 2044 7812
rect 2015 7803 2044 7809
rect 2015 7769 2027 7803
rect 2015 7763 2044 7769
rect 2038 7760 2044 7763
rect 2096 7760 2102 7812
rect 2133 7803 2191 7809
rect 2133 7769 2145 7803
rect 2179 7769 2191 7803
rect 3252 7800 3280 7831
rect 3326 7828 3332 7880
rect 3384 7868 3390 7880
rect 3789 7871 3847 7877
rect 3789 7868 3801 7871
rect 3384 7840 3801 7868
rect 3384 7828 3390 7840
rect 3789 7837 3801 7840
rect 3835 7868 3847 7871
rect 4264 7868 4292 7908
rect 4614 7896 4620 7908
rect 4672 7896 4678 7948
rect 9030 7896 9036 7948
rect 9088 7896 9094 7948
rect 9306 7936 9312 7948
rect 9156 7908 9312 7936
rect 3835 7840 4292 7868
rect 3835 7837 3847 7840
rect 3789 7831 3847 7837
rect 4338 7828 4344 7880
rect 4396 7868 4402 7880
rect 4396 7840 4844 7868
rect 4396 7828 4402 7840
rect 4246 7800 4252 7812
rect 3252 7772 4252 7800
rect 2133 7763 2191 7769
rect 1820 7704 1900 7732
rect 2148 7732 2176 7763
rect 4246 7760 4252 7772
rect 4304 7800 4310 7812
rect 4816 7809 4844 7840
rect 4890 7828 4896 7880
rect 4948 7828 4954 7880
rect 6822 7828 6828 7880
rect 6880 7828 6886 7880
rect 6917 7871 6975 7877
rect 6917 7837 6929 7871
rect 6963 7837 6975 7871
rect 6917 7831 6975 7837
rect 4585 7803 4643 7809
rect 4585 7800 4597 7803
rect 4304 7772 4597 7800
rect 4304 7760 4310 7772
rect 4585 7769 4597 7772
rect 4631 7769 4643 7803
rect 4585 7763 4643 7769
rect 4801 7803 4859 7809
rect 4801 7769 4813 7803
rect 4847 7769 4859 7803
rect 6932 7800 6960 7831
rect 7006 7828 7012 7880
rect 7064 7868 7070 7880
rect 7101 7871 7159 7877
rect 7101 7868 7113 7871
rect 7064 7840 7113 7868
rect 7064 7828 7070 7840
rect 7101 7837 7113 7840
rect 7147 7837 7159 7871
rect 7101 7831 7159 7837
rect 7190 7828 7196 7880
rect 7248 7868 7254 7880
rect 7466 7868 7472 7880
rect 7248 7840 7472 7868
rect 7248 7828 7254 7840
rect 7466 7828 7472 7840
rect 7524 7828 7530 7880
rect 8297 7871 8355 7877
rect 8297 7837 8309 7871
rect 8343 7868 8355 7871
rect 8343 7840 8892 7868
rect 8343 7837 8355 7840
rect 8297 7831 8355 7837
rect 7208 7800 7236 7828
rect 6932 7772 7236 7800
rect 4801 7763 4859 7769
rect 2590 7732 2596 7744
rect 2148 7704 2596 7732
rect 1820 7692 1826 7704
rect 2590 7692 2596 7704
rect 2648 7692 2654 7744
rect 2866 7692 2872 7744
rect 2924 7732 2930 7744
rect 3602 7732 3608 7744
rect 2924 7704 3608 7732
rect 2924 7692 2930 7704
rect 3602 7692 3608 7704
rect 3660 7692 3666 7744
rect 3970 7692 3976 7744
rect 4028 7692 4034 7744
rect 4338 7692 4344 7744
rect 4396 7732 4402 7744
rect 4433 7735 4491 7741
rect 4433 7732 4445 7735
rect 4396 7704 4445 7732
rect 4396 7692 4402 7704
rect 4433 7701 4445 7704
rect 4479 7701 4491 7735
rect 4816 7732 4844 7763
rect 7282 7760 7288 7812
rect 7340 7760 7346 7812
rect 7377 7803 7435 7809
rect 7377 7769 7389 7803
rect 7423 7800 7435 7803
rect 8312 7800 8340 7831
rect 7423 7772 8340 7800
rect 8757 7803 8815 7809
rect 7423 7769 7435 7772
rect 7377 7763 7435 7769
rect 8757 7769 8769 7803
rect 8803 7769 8815 7803
rect 8864 7800 8892 7840
rect 8938 7828 8944 7880
rect 8996 7828 9002 7880
rect 9156 7868 9184 7908
rect 9306 7896 9312 7908
rect 9364 7896 9370 7948
rect 9674 7896 9680 7948
rect 9732 7896 9738 7948
rect 9048 7840 9184 7868
rect 9217 7871 9275 7877
rect 9048 7800 9076 7840
rect 9217 7837 9229 7871
rect 9263 7837 9275 7871
rect 9324 7868 9352 7896
rect 9769 7871 9827 7877
rect 9769 7868 9781 7871
rect 9324 7840 9781 7868
rect 9217 7831 9275 7837
rect 9769 7837 9781 7840
rect 9815 7837 9827 7871
rect 9769 7831 9827 7837
rect 8864 7772 9076 7800
rect 8757 7763 8815 7769
rect 7392 7732 7420 7763
rect 4816 7704 7420 7732
rect 7653 7735 7711 7741
rect 4433 7695 4491 7701
rect 7653 7701 7665 7735
rect 7699 7732 7711 7735
rect 8018 7732 8024 7744
rect 7699 7704 8024 7732
rect 7699 7701 7711 7704
rect 7653 7695 7711 7701
rect 8018 7692 8024 7704
rect 8076 7692 8082 7744
rect 8113 7735 8171 7741
rect 8113 7701 8125 7735
rect 8159 7732 8171 7735
rect 8386 7732 8392 7744
rect 8159 7704 8392 7732
rect 8159 7701 8171 7704
rect 8113 7695 8171 7701
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 8570 7741 8576 7744
rect 8557 7735 8576 7741
rect 8557 7701 8569 7735
rect 8557 7695 8576 7701
rect 8570 7692 8576 7695
rect 8628 7692 8634 7744
rect 8662 7692 8668 7744
rect 8720 7732 8726 7744
rect 8772 7732 8800 7763
rect 9122 7760 9128 7812
rect 9180 7760 9186 7812
rect 9232 7800 9260 7831
rect 12066 7828 12072 7880
rect 12124 7828 12130 7880
rect 12345 7871 12403 7877
rect 12345 7837 12357 7871
rect 12391 7868 12403 7871
rect 12434 7868 12440 7880
rect 12391 7840 12440 7868
rect 12391 7837 12403 7840
rect 12345 7831 12403 7837
rect 12434 7828 12440 7840
rect 12492 7828 12498 7880
rect 12728 7877 12756 7976
rect 13725 7973 13737 8007
rect 13771 7973 13783 8007
rect 13725 7967 13783 7973
rect 12805 7939 12863 7945
rect 12805 7905 12817 7939
rect 12851 7936 12863 7939
rect 13170 7936 13176 7948
rect 12851 7908 13176 7936
rect 12851 7905 12863 7908
rect 12805 7899 12863 7905
rect 13170 7896 13176 7908
rect 13228 7936 13234 7948
rect 13265 7939 13323 7945
rect 13265 7936 13277 7939
rect 13228 7908 13277 7936
rect 13228 7896 13234 7908
rect 13265 7905 13277 7908
rect 13311 7905 13323 7939
rect 13740 7936 13768 7967
rect 14366 7936 14372 7948
rect 13740 7908 14372 7936
rect 13265 7899 13323 7905
rect 14366 7896 14372 7908
rect 14424 7896 14430 7948
rect 14936 7936 14964 8032
rect 15197 7939 15255 7945
rect 15197 7936 15209 7939
rect 14936 7908 15209 7936
rect 15197 7905 15209 7908
rect 15243 7905 15255 7939
rect 15197 7899 15255 7905
rect 15657 7939 15715 7945
rect 15657 7905 15669 7939
rect 15703 7936 15715 7939
rect 15703 7908 15792 7936
rect 15703 7905 15715 7908
rect 15657 7899 15715 7905
rect 12713 7871 12771 7877
rect 12713 7837 12725 7871
rect 12759 7837 12771 7871
rect 12713 7831 12771 7837
rect 12894 7828 12900 7880
rect 12952 7828 12958 7880
rect 13354 7828 13360 7880
rect 13412 7828 13418 7880
rect 13814 7828 13820 7880
rect 13872 7868 13878 7880
rect 14458 7868 14464 7880
rect 13872 7840 14464 7868
rect 13872 7828 13878 7840
rect 14458 7828 14464 7840
rect 14516 7828 14522 7880
rect 14734 7828 14740 7880
rect 14792 7868 14798 7880
rect 15764 7877 15792 7908
rect 15289 7871 15347 7877
rect 15289 7868 15301 7871
rect 14792 7840 15301 7868
rect 14792 7828 14798 7840
rect 15289 7837 15301 7840
rect 15335 7837 15347 7871
rect 15289 7831 15347 7837
rect 15749 7871 15807 7877
rect 15749 7837 15761 7871
rect 15795 7837 15807 7871
rect 15749 7831 15807 7837
rect 9861 7803 9919 7809
rect 9861 7800 9873 7803
rect 9232 7772 9873 7800
rect 9861 7769 9873 7772
rect 9907 7769 9919 7803
rect 9861 7763 9919 7769
rect 9140 7732 9168 7760
rect 8720 7704 9168 7732
rect 8720 7692 8726 7704
rect 12158 7692 12164 7744
rect 12216 7692 12222 7744
rect 15930 7692 15936 7744
rect 15988 7692 15994 7744
rect 1104 7642 16376 7664
rect 1104 7590 3519 7642
rect 3571 7590 3583 7642
rect 3635 7590 3647 7642
rect 3699 7590 3711 7642
rect 3763 7590 3775 7642
rect 3827 7590 7337 7642
rect 7389 7590 7401 7642
rect 7453 7590 7465 7642
rect 7517 7590 7529 7642
rect 7581 7590 7593 7642
rect 7645 7590 11155 7642
rect 11207 7590 11219 7642
rect 11271 7590 11283 7642
rect 11335 7590 11347 7642
rect 11399 7590 11411 7642
rect 11463 7590 14973 7642
rect 15025 7590 15037 7642
rect 15089 7590 15101 7642
rect 15153 7590 15165 7642
rect 15217 7590 15229 7642
rect 15281 7590 16376 7642
rect 1104 7568 16376 7590
rect 2038 7488 2044 7540
rect 2096 7488 2102 7540
rect 2130 7488 2136 7540
rect 2188 7528 2194 7540
rect 2317 7531 2375 7537
rect 2317 7528 2329 7531
rect 2188 7500 2329 7528
rect 2188 7488 2194 7500
rect 2317 7497 2329 7500
rect 2363 7497 2375 7531
rect 2317 7491 2375 7497
rect 2406 7488 2412 7540
rect 2464 7488 2470 7540
rect 3697 7531 3755 7537
rect 3697 7528 3709 7531
rect 2746 7500 3709 7528
rect 934 7420 940 7472
rect 992 7460 998 7472
rect 1489 7463 1547 7469
rect 1489 7460 1501 7463
rect 992 7432 1501 7460
rect 992 7420 998 7432
rect 1489 7429 1501 7432
rect 1535 7429 1547 7463
rect 1489 7423 1547 7429
rect 1854 7420 1860 7472
rect 1912 7420 1918 7472
rect 1946 7420 1952 7472
rect 2004 7420 2010 7472
rect 2056 7460 2084 7488
rect 2746 7460 2774 7500
rect 3697 7497 3709 7500
rect 3743 7497 3755 7531
rect 3697 7491 3755 7497
rect 3878 7488 3884 7540
rect 3936 7488 3942 7540
rect 3970 7488 3976 7540
rect 4028 7488 4034 7540
rect 4154 7488 4160 7540
rect 4212 7528 4218 7540
rect 4525 7531 4583 7537
rect 4525 7528 4537 7531
rect 4212 7500 4537 7528
rect 4212 7488 4218 7500
rect 4525 7497 4537 7500
rect 4571 7497 4583 7531
rect 4525 7491 4583 7497
rect 4890 7488 4896 7540
rect 4948 7488 4954 7540
rect 5534 7488 5540 7540
rect 5592 7528 5598 7540
rect 5592 7500 5672 7528
rect 5592 7488 5598 7500
rect 2056 7432 2774 7460
rect 2866 7420 2872 7472
rect 2924 7420 2930 7472
rect 3085 7463 3143 7469
rect 3085 7429 3097 7463
rect 3131 7460 3143 7463
rect 3131 7432 3832 7460
rect 3131 7429 3143 7432
rect 3085 7423 3143 7429
rect 1762 7352 1768 7404
rect 1820 7352 1826 7404
rect 1872 7392 1900 7420
rect 3804 7404 3832 7432
rect 2041 7395 2099 7401
rect 2041 7392 2053 7395
rect 1872 7364 2053 7392
rect 2041 7361 2053 7364
rect 2087 7361 2099 7395
rect 2041 7355 2099 7361
rect 2133 7395 2191 7401
rect 2133 7361 2145 7395
rect 2179 7392 2191 7395
rect 2409 7395 2467 7401
rect 2409 7392 2421 7395
rect 2179 7364 2421 7392
rect 2179 7361 2191 7364
rect 2133 7355 2191 7361
rect 2409 7361 2421 7364
rect 2455 7392 2467 7395
rect 2498 7392 2504 7404
rect 2455 7364 2504 7392
rect 2455 7361 2467 7364
rect 2409 7355 2467 7361
rect 2498 7352 2504 7364
rect 2556 7352 2562 7404
rect 2593 7395 2651 7401
rect 2593 7361 2605 7395
rect 2639 7392 2651 7395
rect 2639 7364 3464 7392
rect 2639 7361 2651 7364
rect 2593 7355 2651 7361
rect 1673 7327 1731 7333
rect 1673 7293 1685 7327
rect 1719 7324 1731 7327
rect 2314 7324 2320 7336
rect 1719 7296 2320 7324
rect 1719 7293 1731 7296
rect 1673 7287 1731 7293
rect 2314 7284 2320 7296
rect 2372 7324 2378 7336
rect 2608 7324 2636 7355
rect 2372 7296 2636 7324
rect 2372 7284 2378 7296
rect 3237 7259 3295 7265
rect 3237 7225 3249 7259
rect 3283 7256 3295 7259
rect 3326 7256 3332 7268
rect 3283 7228 3332 7256
rect 3283 7225 3295 7228
rect 3237 7219 3295 7225
rect 3326 7216 3332 7228
rect 3384 7216 3390 7268
rect 3436 7256 3464 7364
rect 3786 7352 3792 7404
rect 3844 7352 3850 7404
rect 3896 7401 3924 7488
rect 3988 7460 4016 7488
rect 4908 7460 4936 7488
rect 5644 7469 5672 7500
rect 5902 7488 5908 7540
rect 5960 7528 5966 7540
rect 6089 7531 6147 7537
rect 6089 7528 6101 7531
rect 5960 7500 6101 7528
rect 5960 7488 5966 7500
rect 6089 7497 6101 7500
rect 6135 7528 6147 7531
rect 6454 7528 6460 7540
rect 6135 7500 6460 7528
rect 6135 7497 6147 7500
rect 6089 7491 6147 7497
rect 6454 7488 6460 7500
rect 6512 7488 6518 7540
rect 7558 7488 7564 7540
rect 7616 7488 7622 7540
rect 8754 7528 8760 7540
rect 7668 7500 8760 7528
rect 3988 7432 4476 7460
rect 4448 7401 4476 7432
rect 4816 7432 4936 7460
rect 5629 7463 5687 7469
rect 3889 7395 3947 7401
rect 3889 7361 3901 7395
rect 3935 7361 3947 7395
rect 3889 7355 3947 7361
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7392 4215 7395
rect 4433 7395 4491 7401
rect 4203 7364 4292 7392
rect 4203 7361 4215 7364
rect 4157 7355 4215 7361
rect 4264 7336 4292 7364
rect 4433 7361 4445 7395
rect 4479 7361 4491 7395
rect 4433 7355 4491 7361
rect 4522 7352 4528 7404
rect 4580 7392 4586 7404
rect 4617 7395 4675 7401
rect 4617 7392 4629 7395
rect 4580 7364 4629 7392
rect 4580 7352 4586 7364
rect 4617 7361 4629 7364
rect 4663 7361 4675 7395
rect 4617 7355 4675 7361
rect 4709 7395 4767 7401
rect 4709 7361 4721 7395
rect 4755 7392 4767 7395
rect 4816 7392 4844 7432
rect 5629 7429 5641 7463
rect 5675 7429 5687 7463
rect 5629 7423 5687 7429
rect 5721 7463 5779 7469
rect 5721 7429 5733 7463
rect 5767 7460 5779 7463
rect 7469 7463 7527 7469
rect 5767 7432 6592 7460
rect 5767 7429 5779 7432
rect 5721 7423 5779 7429
rect 4755 7364 4844 7392
rect 4893 7395 4951 7401
rect 4755 7361 4767 7364
rect 4709 7355 4767 7361
rect 4893 7361 4905 7395
rect 4939 7361 4951 7395
rect 4893 7355 4951 7361
rect 3970 7284 3976 7336
rect 4028 7284 4034 7336
rect 4246 7284 4252 7336
rect 4304 7284 4310 7336
rect 4724 7256 4752 7355
rect 4908 7324 4936 7355
rect 5442 7352 5448 7404
rect 5500 7392 5506 7404
rect 5537 7395 5595 7401
rect 5537 7392 5549 7395
rect 5500 7364 5549 7392
rect 5500 7352 5506 7364
rect 5537 7361 5549 7364
rect 5583 7361 5595 7395
rect 5537 7355 5595 7361
rect 5810 7352 5816 7404
rect 5868 7392 5874 7404
rect 5905 7395 5963 7401
rect 5905 7392 5917 7395
rect 5868 7364 5917 7392
rect 5868 7352 5874 7364
rect 5905 7361 5917 7364
rect 5951 7361 5963 7395
rect 5905 7355 5963 7361
rect 5997 7395 6055 7401
rect 5997 7361 6009 7395
rect 6043 7392 6055 7395
rect 6365 7395 6423 7401
rect 6365 7392 6377 7395
rect 6043 7364 6377 7392
rect 6043 7361 6055 7364
rect 5997 7355 6055 7361
rect 6365 7361 6377 7364
rect 6411 7361 6423 7395
rect 6365 7355 6423 7361
rect 6012 7324 6040 7355
rect 4908 7296 6040 7324
rect 3436 7228 4752 7256
rect 5644 7200 5672 7296
rect 6564 7200 6592 7432
rect 7469 7429 7481 7463
rect 7515 7460 7527 7463
rect 7576 7460 7604 7488
rect 7515 7432 7604 7460
rect 7515 7429 7527 7432
rect 7469 7423 7527 7429
rect 7668 7423 7696 7500
rect 8754 7488 8760 7500
rect 8812 7528 8818 7540
rect 9030 7528 9036 7540
rect 8812 7500 9036 7528
rect 8812 7488 8818 7500
rect 9030 7488 9036 7500
rect 9088 7488 9094 7540
rect 9861 7531 9919 7537
rect 9861 7497 9873 7531
rect 9907 7528 9919 7531
rect 10042 7528 10048 7540
rect 9907 7500 10048 7528
rect 9907 7497 9919 7500
rect 9861 7491 9919 7497
rect 10042 7488 10048 7500
rect 10100 7528 10106 7540
rect 10100 7500 10364 7528
rect 10100 7488 10106 7500
rect 7658 7417 7716 7423
rect 8018 7420 8024 7472
rect 8076 7420 8082 7472
rect 8294 7420 8300 7472
rect 8352 7460 8358 7472
rect 8478 7460 8484 7472
rect 8352 7432 8484 7460
rect 8352 7420 8358 7432
rect 8478 7420 8484 7432
rect 8536 7460 8542 7472
rect 8849 7463 8907 7469
rect 8849 7460 8861 7463
rect 8536 7432 8861 7460
rect 8536 7420 8542 7432
rect 8849 7429 8861 7432
rect 8895 7429 8907 7463
rect 9490 7460 9496 7472
rect 8849 7423 8907 7429
rect 8956 7432 9496 7460
rect 7282 7352 7288 7404
rect 7340 7352 7346 7404
rect 7558 7352 7564 7404
rect 7616 7352 7622 7404
rect 7658 7383 7670 7417
rect 7704 7383 7716 7417
rect 7658 7377 7716 7383
rect 8036 7392 8064 7420
rect 8956 7392 8984 7432
rect 9490 7420 9496 7432
rect 9548 7420 9554 7472
rect 10336 7469 10364 7500
rect 12434 7488 12440 7540
rect 12492 7537 12498 7540
rect 12492 7531 12511 7537
rect 12499 7497 12511 7531
rect 12492 7491 12511 7497
rect 12621 7531 12679 7537
rect 12621 7497 12633 7531
rect 12667 7528 12679 7531
rect 12894 7528 12900 7540
rect 12667 7500 12900 7528
rect 12667 7497 12679 7500
rect 12621 7491 12679 7497
rect 12492 7488 12498 7491
rect 12894 7488 12900 7500
rect 12952 7488 12958 7540
rect 13170 7488 13176 7540
rect 13228 7488 13234 7540
rect 13630 7488 13636 7540
rect 13688 7488 13694 7540
rect 14366 7488 14372 7540
rect 14424 7488 14430 7540
rect 14826 7488 14832 7540
rect 14884 7528 14890 7540
rect 14921 7531 14979 7537
rect 14921 7528 14933 7531
rect 14884 7500 14933 7528
rect 14884 7488 14890 7500
rect 14921 7497 14933 7500
rect 14967 7497 14979 7531
rect 14921 7491 14979 7497
rect 9693 7463 9751 7469
rect 9693 7460 9705 7463
rect 9600 7432 9705 7460
rect 8036 7364 8984 7392
rect 9033 7395 9091 7401
rect 9033 7361 9045 7395
rect 9079 7361 9091 7395
rect 9033 7355 9091 7361
rect 7377 7327 7435 7333
rect 7377 7293 7389 7327
rect 7423 7324 7435 7327
rect 9048 7324 9076 7355
rect 9306 7352 9312 7404
rect 9364 7392 9370 7404
rect 9600 7392 9628 7432
rect 9693 7429 9705 7432
rect 9739 7429 9751 7463
rect 9693 7423 9751 7429
rect 10321 7463 10379 7469
rect 10321 7429 10333 7463
rect 10367 7429 10379 7463
rect 10870 7460 10876 7472
rect 10321 7423 10379 7429
rect 10428 7432 10876 7460
rect 9364 7364 9628 7392
rect 9364 7352 9370 7364
rect 10134 7352 10140 7404
rect 10192 7352 10198 7404
rect 7423 7296 9076 7324
rect 9217 7327 9275 7333
rect 7423 7293 7435 7296
rect 7377 7287 7435 7293
rect 9217 7293 9229 7327
rect 9263 7324 9275 7327
rect 10428 7324 10456 7432
rect 10870 7420 10876 7432
rect 10928 7460 10934 7472
rect 11149 7463 11207 7469
rect 11149 7460 11161 7463
rect 10928 7432 11161 7460
rect 10928 7420 10934 7432
rect 11149 7429 11161 7432
rect 11195 7429 11207 7463
rect 11149 7423 11207 7429
rect 11333 7463 11391 7469
rect 11333 7429 11345 7463
rect 11379 7460 11391 7463
rect 12158 7460 12164 7472
rect 11379 7432 12164 7460
rect 11379 7429 11391 7432
rect 11333 7423 11391 7429
rect 12158 7420 12164 7432
rect 12216 7460 12222 7472
rect 12253 7463 12311 7469
rect 12253 7460 12265 7463
rect 12216 7432 12265 7460
rect 12216 7420 12222 7432
rect 12253 7429 12265 7432
rect 12299 7429 12311 7463
rect 12253 7423 12311 7429
rect 13188 7401 13216 7488
rect 10965 7395 11023 7401
rect 10965 7392 10977 7395
rect 9263 7296 10456 7324
rect 10520 7364 10977 7392
rect 9263 7293 9275 7296
rect 9217 7287 9275 7293
rect 7006 7216 7012 7268
rect 7064 7256 7070 7268
rect 7834 7256 7840 7268
rect 7064 7228 7840 7256
rect 7064 7216 7070 7228
rect 7834 7216 7840 7228
rect 7892 7216 7898 7268
rect 2774 7148 2780 7200
rect 2832 7188 2838 7200
rect 3053 7191 3111 7197
rect 3053 7188 3065 7191
rect 2832 7160 3065 7188
rect 2832 7148 2838 7160
rect 3053 7157 3065 7160
rect 3099 7157 3111 7191
rect 3053 7151 3111 7157
rect 3786 7148 3792 7200
rect 3844 7188 3850 7200
rect 4062 7188 4068 7200
rect 3844 7160 4068 7188
rect 3844 7148 3850 7160
rect 4062 7148 4068 7160
rect 4120 7188 4126 7200
rect 4341 7191 4399 7197
rect 4341 7188 4353 7191
rect 4120 7160 4353 7188
rect 4120 7148 4126 7160
rect 4341 7157 4353 7160
rect 4387 7188 4399 7191
rect 4706 7188 4712 7200
rect 4387 7160 4712 7188
rect 4387 7157 4399 7160
rect 4341 7151 4399 7157
rect 4706 7148 4712 7160
rect 4764 7148 4770 7200
rect 4798 7148 4804 7200
rect 4856 7148 4862 7200
rect 4890 7148 4896 7200
rect 4948 7188 4954 7200
rect 5353 7191 5411 7197
rect 5353 7188 5365 7191
rect 4948 7160 5365 7188
rect 4948 7148 4954 7160
rect 5353 7157 5365 7160
rect 5399 7157 5411 7191
rect 5353 7151 5411 7157
rect 5626 7148 5632 7200
rect 5684 7148 5690 7200
rect 5810 7148 5816 7200
rect 5868 7188 5874 7200
rect 6178 7188 6184 7200
rect 5868 7160 6184 7188
rect 5868 7148 5874 7160
rect 6178 7148 6184 7160
rect 6236 7148 6242 7200
rect 6546 7148 6552 7200
rect 6604 7188 6610 7200
rect 7282 7188 7288 7200
rect 6604 7160 7288 7188
rect 6604 7148 6610 7160
rect 7282 7148 7288 7160
rect 7340 7188 7346 7200
rect 8662 7188 8668 7200
rect 7340 7160 8668 7188
rect 7340 7148 7346 7160
rect 8662 7148 8668 7160
rect 8720 7148 8726 7200
rect 9674 7148 9680 7200
rect 9732 7148 9738 7200
rect 10410 7148 10416 7200
rect 10468 7188 10474 7200
rect 10520 7197 10548 7364
rect 10965 7361 10977 7364
rect 11011 7361 11023 7395
rect 10965 7355 11023 7361
rect 13173 7395 13231 7401
rect 13173 7361 13185 7395
rect 13219 7361 13231 7395
rect 13173 7355 13231 7361
rect 12802 7216 12808 7268
rect 12860 7256 12866 7268
rect 13354 7256 13360 7268
rect 12860 7228 13360 7256
rect 12860 7216 12866 7228
rect 13354 7216 13360 7228
rect 13412 7256 13418 7268
rect 13449 7259 13507 7265
rect 13449 7256 13461 7259
rect 13412 7228 13461 7256
rect 13412 7216 13418 7228
rect 13449 7225 13461 7228
rect 13495 7225 13507 7259
rect 14384 7256 14412 7488
rect 14458 7420 14464 7472
rect 14516 7420 14522 7472
rect 14737 7259 14795 7265
rect 14737 7256 14749 7259
rect 14384 7228 14749 7256
rect 13449 7219 13507 7225
rect 14737 7225 14749 7228
rect 14783 7225 14795 7259
rect 14737 7219 14795 7225
rect 10505 7191 10563 7197
rect 10505 7188 10517 7191
rect 10468 7160 10517 7188
rect 10468 7148 10474 7160
rect 10505 7157 10517 7160
rect 10551 7157 10563 7191
rect 10505 7151 10563 7157
rect 12066 7148 12072 7200
rect 12124 7188 12130 7200
rect 12437 7191 12495 7197
rect 12437 7188 12449 7191
rect 12124 7160 12449 7188
rect 12124 7148 12130 7160
rect 12437 7157 12449 7160
rect 12483 7157 12495 7191
rect 12437 7151 12495 7157
rect 1104 7098 16376 7120
rect 1104 7046 2859 7098
rect 2911 7046 2923 7098
rect 2975 7046 2987 7098
rect 3039 7046 3051 7098
rect 3103 7046 3115 7098
rect 3167 7046 6677 7098
rect 6729 7046 6741 7098
rect 6793 7046 6805 7098
rect 6857 7046 6869 7098
rect 6921 7046 6933 7098
rect 6985 7046 10495 7098
rect 10547 7046 10559 7098
rect 10611 7046 10623 7098
rect 10675 7046 10687 7098
rect 10739 7046 10751 7098
rect 10803 7046 14313 7098
rect 14365 7046 14377 7098
rect 14429 7046 14441 7098
rect 14493 7046 14505 7098
rect 14557 7046 14569 7098
rect 14621 7046 16376 7098
rect 1104 7024 16376 7046
rect 1854 6944 1860 6996
rect 1912 6984 1918 6996
rect 3326 6984 3332 6996
rect 1912 6956 3332 6984
rect 1912 6944 1918 6956
rect 3326 6944 3332 6956
rect 3384 6984 3390 6996
rect 3970 6984 3976 6996
rect 3384 6956 3976 6984
rect 3384 6944 3390 6956
rect 3970 6944 3976 6956
rect 4028 6984 4034 6996
rect 5810 6984 5816 6996
rect 4028 6956 5816 6984
rect 4028 6944 4034 6956
rect 5810 6944 5816 6956
rect 5868 6944 5874 6996
rect 6086 6944 6092 6996
rect 6144 6944 6150 6996
rect 6178 6944 6184 6996
rect 6236 6984 6242 6996
rect 7742 6984 7748 6996
rect 6236 6956 7748 6984
rect 6236 6944 6242 6956
rect 7742 6944 7748 6956
rect 7800 6944 7806 6996
rect 9309 6987 9367 6993
rect 9309 6953 9321 6987
rect 9355 6984 9367 6987
rect 10134 6984 10140 6996
rect 9355 6956 10140 6984
rect 9355 6953 9367 6956
rect 9309 6947 9367 6953
rect 10134 6944 10140 6956
rect 10192 6944 10198 6996
rect 12066 6944 12072 6996
rect 12124 6984 12130 6996
rect 12161 6987 12219 6993
rect 12161 6984 12173 6987
rect 12124 6956 12173 6984
rect 12124 6944 12130 6956
rect 12161 6953 12173 6956
rect 12207 6953 12219 6987
rect 12161 6947 12219 6953
rect 2682 6876 2688 6928
rect 2740 6916 2746 6928
rect 3053 6919 3111 6925
rect 3053 6916 3065 6919
rect 2740 6888 3065 6916
rect 2740 6876 2746 6888
rect 3053 6885 3065 6888
rect 3099 6885 3111 6919
rect 3053 6879 3111 6885
rect 4172 6888 4660 6916
rect 1762 6808 1768 6860
rect 1820 6848 1826 6860
rect 2038 6848 2044 6860
rect 1820 6820 2044 6848
rect 1820 6808 1826 6820
rect 2038 6808 2044 6820
rect 2096 6808 2102 6860
rect 4172 6848 4200 6888
rect 3068 6820 3280 6848
rect 1854 6740 1860 6792
rect 1912 6780 1918 6792
rect 2225 6783 2283 6789
rect 2225 6780 2237 6783
rect 1912 6752 2237 6780
rect 1912 6740 1918 6752
rect 2225 6749 2237 6752
rect 2271 6780 2283 6783
rect 2961 6783 3019 6789
rect 2961 6780 2973 6783
rect 2271 6752 2973 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 2961 6749 2973 6752
rect 3007 6749 3019 6783
rect 2961 6743 3019 6749
rect 1762 6672 1768 6724
rect 1820 6712 1826 6724
rect 2501 6715 2559 6721
rect 2501 6712 2513 6715
rect 1820 6684 2513 6712
rect 1820 6672 1826 6684
rect 2501 6681 2513 6684
rect 2547 6712 2559 6715
rect 3068 6712 3096 6820
rect 3252 6789 3280 6820
rect 3988 6820 4200 6848
rect 3988 6792 4016 6820
rect 3136 6783 3194 6789
rect 3136 6749 3148 6783
rect 3182 6749 3194 6783
rect 3136 6743 3194 6749
rect 3237 6783 3295 6789
rect 3237 6749 3249 6783
rect 3283 6749 3295 6783
rect 3237 6743 3295 6749
rect 2547 6684 3096 6712
rect 3160 6712 3188 6743
rect 3878 6740 3884 6792
rect 3936 6740 3942 6792
rect 3970 6740 3976 6792
rect 4028 6740 4034 6792
rect 4154 6740 4160 6792
rect 4212 6740 4218 6792
rect 4430 6740 4436 6792
rect 4488 6780 4494 6792
rect 4632 6789 4660 6888
rect 5534 6876 5540 6928
rect 5592 6916 5598 6928
rect 6454 6916 6460 6928
rect 5592 6888 6460 6916
rect 5592 6876 5598 6888
rect 6454 6876 6460 6888
rect 6512 6916 6518 6928
rect 7558 6916 7564 6928
rect 6512 6888 7564 6916
rect 6512 6876 6518 6888
rect 7558 6876 7564 6888
rect 7616 6916 7622 6928
rect 8110 6916 8116 6928
rect 7616 6888 8116 6916
rect 7616 6876 7622 6888
rect 8110 6876 8116 6888
rect 8168 6876 8174 6928
rect 9674 6916 9680 6928
rect 9600 6888 9680 6916
rect 4706 6808 4712 6860
rect 4764 6848 4770 6860
rect 6362 6848 6368 6860
rect 4764 6820 5212 6848
rect 4764 6808 4770 6820
rect 4525 6783 4583 6789
rect 4525 6780 4537 6783
rect 4488 6752 4537 6780
rect 4488 6740 4494 6752
rect 4525 6749 4537 6752
rect 4571 6749 4583 6783
rect 4525 6743 4583 6749
rect 4617 6783 4675 6789
rect 4617 6749 4629 6783
rect 4663 6749 4675 6783
rect 4617 6743 4675 6749
rect 4798 6740 4804 6792
rect 4856 6780 4862 6792
rect 5184 6789 5212 6820
rect 5276 6820 6368 6848
rect 4985 6783 5043 6789
rect 4985 6780 4997 6783
rect 4856 6752 4997 6780
rect 4856 6740 4862 6752
rect 4985 6749 4997 6752
rect 5031 6749 5043 6783
rect 4985 6743 5043 6749
rect 5169 6783 5227 6789
rect 5169 6749 5181 6783
rect 5215 6749 5227 6783
rect 5169 6743 5227 6749
rect 3896 6712 3924 6740
rect 5276 6712 5304 6820
rect 5350 6740 5356 6792
rect 5408 6780 5414 6792
rect 5445 6783 5503 6789
rect 5445 6780 5457 6783
rect 5408 6752 5457 6780
rect 5408 6740 5414 6752
rect 5445 6749 5457 6752
rect 5491 6749 5503 6783
rect 5445 6743 5503 6749
rect 5534 6740 5540 6792
rect 5592 6740 5598 6792
rect 5828 6789 5856 6820
rect 6362 6808 6368 6820
rect 6420 6808 6426 6860
rect 6914 6857 6920 6860
rect 6897 6851 6920 6857
rect 6897 6817 6909 6851
rect 6897 6811 6920 6817
rect 6914 6808 6920 6811
rect 6972 6808 6978 6860
rect 8021 6851 8079 6857
rect 8021 6817 8033 6851
rect 8067 6848 8079 6851
rect 8067 6820 8248 6848
rect 8067 6817 8079 6820
rect 8021 6811 8079 6817
rect 5813 6783 5871 6789
rect 5813 6749 5825 6783
rect 5859 6780 5871 6783
rect 5905 6783 5963 6789
rect 5905 6780 5917 6783
rect 5859 6752 5917 6780
rect 5859 6749 5871 6752
rect 5813 6743 5871 6749
rect 5905 6749 5917 6752
rect 5951 6749 5963 6783
rect 7101 6783 7159 6789
rect 7101 6780 7113 6783
rect 5905 6743 5963 6749
rect 6012 6752 7113 6780
rect 3160 6684 3280 6712
rect 3896 6684 5304 6712
rect 2547 6681 2559 6684
rect 2501 6675 2559 6681
rect 3252 6656 3280 6684
rect 5626 6672 5632 6724
rect 5684 6672 5690 6724
rect 2682 6604 2688 6656
rect 2740 6644 2746 6656
rect 2777 6647 2835 6653
rect 2777 6644 2789 6647
rect 2740 6616 2789 6644
rect 2740 6604 2746 6616
rect 2777 6613 2789 6616
rect 2823 6613 2835 6647
rect 2777 6607 2835 6613
rect 3234 6604 3240 6656
rect 3292 6604 3298 6656
rect 3329 6647 3387 6653
rect 3329 6613 3341 6647
rect 3375 6644 3387 6647
rect 4522 6644 4528 6656
rect 3375 6616 4528 6644
rect 3375 6613 3387 6616
rect 3329 6607 3387 6613
rect 4522 6604 4528 6616
rect 4580 6604 4586 6656
rect 5074 6604 5080 6656
rect 5132 6604 5138 6656
rect 5258 6604 5264 6656
rect 5316 6644 5322 6656
rect 6012 6644 6040 6752
rect 7101 6749 7113 6752
rect 7147 6749 7159 6783
rect 7101 6743 7159 6749
rect 7929 6783 7987 6789
rect 7929 6749 7941 6783
rect 7975 6780 7987 6783
rect 7975 6752 8064 6780
rect 7975 6749 7987 6752
rect 7929 6743 7987 6749
rect 6822 6672 6828 6724
rect 6880 6672 6886 6724
rect 8036 6656 8064 6752
rect 8110 6740 8116 6792
rect 8168 6740 8174 6792
rect 8220 6789 8248 6820
rect 8205 6783 8263 6789
rect 8205 6749 8217 6783
rect 8251 6780 8263 6783
rect 8570 6780 8576 6792
rect 8251 6752 8576 6780
rect 8251 6749 8263 6752
rect 8205 6743 8263 6749
rect 8570 6740 8576 6752
rect 8628 6740 8634 6792
rect 9490 6740 9496 6792
rect 9548 6740 9554 6792
rect 9600 6789 9628 6888
rect 9674 6876 9680 6888
rect 9732 6876 9738 6928
rect 9585 6783 9643 6789
rect 9585 6749 9597 6783
rect 9631 6749 9643 6783
rect 9585 6743 9643 6749
rect 10410 6740 10416 6792
rect 10468 6780 10474 6792
rect 10689 6783 10747 6789
rect 10689 6780 10701 6783
rect 10468 6752 10701 6780
rect 10468 6740 10474 6752
rect 10689 6749 10701 6752
rect 10735 6749 10747 6783
rect 10689 6743 10747 6749
rect 10870 6740 10876 6792
rect 10928 6740 10934 6792
rect 11793 6783 11851 6789
rect 11793 6780 11805 6783
rect 11716 6752 11805 6780
rect 8754 6672 8760 6724
rect 8812 6712 8818 6724
rect 9306 6712 9312 6724
rect 8812 6684 9312 6712
rect 8812 6672 8818 6684
rect 9306 6672 9312 6684
rect 9364 6672 9370 6724
rect 5316 6616 6040 6644
rect 5316 6604 5322 6616
rect 7006 6604 7012 6656
rect 7064 6604 7070 6656
rect 8018 6604 8024 6656
rect 8076 6604 8082 6656
rect 8294 6604 8300 6656
rect 8352 6604 8358 6656
rect 11606 6604 11612 6656
rect 11664 6644 11670 6656
rect 11716 6653 11744 6752
rect 11793 6749 11805 6752
rect 11839 6749 11851 6783
rect 11793 6743 11851 6749
rect 11885 6783 11943 6789
rect 11885 6749 11897 6783
rect 11931 6780 11943 6783
rect 12069 6783 12127 6789
rect 12069 6780 12081 6783
rect 11931 6752 12081 6780
rect 11931 6749 11943 6752
rect 11885 6743 11943 6749
rect 12069 6749 12081 6752
rect 12115 6749 12127 6783
rect 12069 6743 12127 6749
rect 12250 6740 12256 6792
rect 12308 6740 12314 6792
rect 11701 6647 11759 6653
rect 11701 6644 11713 6647
rect 11664 6616 11713 6644
rect 11664 6604 11670 6616
rect 11701 6613 11713 6616
rect 11747 6613 11759 6647
rect 11701 6607 11759 6613
rect 1104 6554 16376 6576
rect 1104 6502 3519 6554
rect 3571 6502 3583 6554
rect 3635 6502 3647 6554
rect 3699 6502 3711 6554
rect 3763 6502 3775 6554
rect 3827 6502 7337 6554
rect 7389 6502 7401 6554
rect 7453 6502 7465 6554
rect 7517 6502 7529 6554
rect 7581 6502 7593 6554
rect 7645 6502 11155 6554
rect 11207 6502 11219 6554
rect 11271 6502 11283 6554
rect 11335 6502 11347 6554
rect 11399 6502 11411 6554
rect 11463 6502 14973 6554
rect 15025 6502 15037 6554
rect 15089 6502 15101 6554
rect 15153 6502 15165 6554
rect 15217 6502 15229 6554
rect 15281 6502 16376 6554
rect 1104 6480 16376 6502
rect 2314 6400 2320 6452
rect 2372 6440 2378 6452
rect 2409 6443 2467 6449
rect 2409 6440 2421 6443
rect 2372 6412 2421 6440
rect 2372 6400 2378 6412
rect 2409 6409 2421 6412
rect 2455 6409 2467 6443
rect 4154 6440 4160 6452
rect 2409 6403 2467 6409
rect 2792 6412 4160 6440
rect 934 6264 940 6316
rect 992 6304 998 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 992 6276 1409 6304
rect 992 6264 998 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 1854 6264 1860 6316
rect 1912 6304 1918 6316
rect 2225 6307 2283 6313
rect 2225 6304 2237 6307
rect 1912 6276 2237 6304
rect 1912 6264 1918 6276
rect 2225 6273 2237 6276
rect 2271 6273 2283 6307
rect 2225 6267 2283 6273
rect 2314 6264 2320 6316
rect 2372 6264 2378 6316
rect 2792 6304 2820 6412
rect 4154 6400 4160 6412
rect 4212 6400 4218 6452
rect 4706 6440 4712 6452
rect 4632 6412 4712 6440
rect 3421 6375 3479 6381
rect 3421 6341 3433 6375
rect 3467 6372 3479 6375
rect 3878 6372 3884 6384
rect 3467 6344 3884 6372
rect 3467 6341 3479 6344
rect 3421 6335 3479 6341
rect 3878 6332 3884 6344
rect 3936 6332 3942 6384
rect 4632 6381 4660 6412
rect 4706 6400 4712 6412
rect 4764 6400 4770 6452
rect 5537 6443 5595 6449
rect 5537 6440 5549 6443
rect 4816 6412 5549 6440
rect 4816 6381 4844 6412
rect 5537 6409 5549 6412
rect 5583 6440 5595 6443
rect 7006 6440 7012 6452
rect 5583 6412 7012 6440
rect 5583 6409 5595 6412
rect 5537 6403 5595 6409
rect 7006 6400 7012 6412
rect 7064 6400 7070 6452
rect 7098 6400 7104 6452
rect 7156 6440 7162 6452
rect 7469 6443 7527 6449
rect 7469 6440 7481 6443
rect 7156 6412 7481 6440
rect 7156 6400 7162 6412
rect 7469 6409 7481 6412
rect 7515 6409 7527 6443
rect 7469 6403 7527 6409
rect 7926 6400 7932 6452
rect 7984 6440 7990 6452
rect 8205 6443 8263 6449
rect 8205 6440 8217 6443
rect 7984 6412 8217 6440
rect 7984 6400 7990 6412
rect 8205 6409 8217 6412
rect 8251 6409 8263 6443
rect 8205 6403 8263 6409
rect 8294 6400 8300 6452
rect 8352 6440 8358 6452
rect 8639 6443 8697 6449
rect 8639 6440 8651 6443
rect 8352 6412 8651 6440
rect 8352 6400 8358 6412
rect 8639 6409 8651 6412
rect 8685 6409 8697 6443
rect 8639 6403 8697 6409
rect 9030 6400 9036 6452
rect 9088 6400 9094 6452
rect 12802 6400 12808 6452
rect 12860 6400 12866 6452
rect 14734 6400 14740 6452
rect 14792 6440 14798 6452
rect 14829 6443 14887 6449
rect 14829 6440 14841 6443
rect 14792 6412 14841 6440
rect 14792 6400 14798 6412
rect 14829 6409 14841 6412
rect 14875 6409 14887 6443
rect 14829 6403 14887 6409
rect 4617 6375 4675 6381
rect 4617 6341 4629 6375
rect 4663 6341 4675 6375
rect 4617 6335 4675 6341
rect 4801 6375 4859 6381
rect 4801 6341 4813 6375
rect 4847 6341 4859 6375
rect 4801 6335 4859 6341
rect 4982 6332 4988 6384
rect 5040 6381 5046 6384
rect 5040 6375 5075 6381
rect 5063 6372 5075 6375
rect 6822 6372 6828 6384
rect 5063 6344 6828 6372
rect 5063 6341 5075 6344
rect 5040 6335 5075 6341
rect 5040 6332 5046 6335
rect 6822 6332 6828 6344
rect 6880 6332 6886 6384
rect 8846 6332 8852 6384
rect 8904 6332 8910 6384
rect 10042 6372 10048 6384
rect 9140 6344 10048 6372
rect 2869 6307 2927 6313
rect 2869 6304 2881 6307
rect 2608 6276 2881 6304
rect 1670 6196 1676 6248
rect 1728 6196 1734 6248
rect 1946 6196 1952 6248
rect 2004 6236 2010 6248
rect 2608 6245 2636 6276
rect 2869 6273 2881 6276
rect 2915 6273 2927 6307
rect 3697 6307 3755 6313
rect 3697 6304 3709 6307
rect 2869 6267 2927 6273
rect 3436 6276 3709 6304
rect 2593 6239 2651 6245
rect 2593 6236 2605 6239
rect 2004 6208 2605 6236
rect 2004 6196 2010 6208
rect 2593 6205 2605 6208
rect 2639 6205 2651 6239
rect 2593 6199 2651 6205
rect 2685 6239 2743 6245
rect 2685 6205 2697 6239
rect 2731 6236 2743 6239
rect 3234 6236 3240 6248
rect 2731 6208 3240 6236
rect 2731 6205 2743 6208
rect 2685 6199 2743 6205
rect 3234 6196 3240 6208
rect 3292 6196 3298 6248
rect 3436 6112 3464 6276
rect 3697 6273 3709 6276
rect 3743 6304 3755 6307
rect 3970 6304 3976 6316
rect 3743 6276 3976 6304
rect 3743 6273 3755 6276
rect 3697 6267 3755 6273
rect 3970 6264 3976 6276
rect 4028 6264 4034 6316
rect 4433 6307 4491 6313
rect 4433 6273 4445 6307
rect 4479 6273 4491 6307
rect 4433 6267 4491 6273
rect 3881 6239 3939 6245
rect 3881 6205 3893 6239
rect 3927 6236 3939 6239
rect 4154 6236 4160 6248
rect 3927 6208 4160 6236
rect 3927 6205 3939 6208
rect 3881 6199 3939 6205
rect 4154 6196 4160 6208
rect 4212 6196 4218 6248
rect 4448 6112 4476 6267
rect 4522 6264 4528 6316
rect 4580 6304 4586 6316
rect 5721 6307 5779 6313
rect 5721 6304 5733 6307
rect 4580 6276 5733 6304
rect 4580 6264 4586 6276
rect 5721 6273 5733 6276
rect 5767 6273 5779 6307
rect 5721 6267 5779 6273
rect 5258 6196 5264 6248
rect 5316 6196 5322 6248
rect 5350 6196 5356 6248
rect 5408 6196 5414 6248
rect 5736 6236 5764 6267
rect 5902 6264 5908 6316
rect 5960 6264 5966 6316
rect 5997 6307 6055 6313
rect 5997 6273 6009 6307
rect 6043 6304 6055 6307
rect 6178 6304 6184 6316
rect 6043 6276 6184 6304
rect 6043 6273 6055 6276
rect 5997 6267 6055 6273
rect 6178 6264 6184 6276
rect 6236 6264 6242 6316
rect 6362 6264 6368 6316
rect 6420 6264 6426 6316
rect 6454 6264 6460 6316
rect 6512 6304 6518 6316
rect 6549 6307 6607 6313
rect 6549 6304 6561 6307
rect 6512 6276 6561 6304
rect 6512 6264 6518 6276
rect 6549 6273 6561 6276
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 6638 6264 6644 6316
rect 6696 6264 6702 6316
rect 6730 6264 6736 6316
rect 6788 6264 6794 6316
rect 7834 6264 7840 6316
rect 7892 6264 7898 6316
rect 8018 6264 8024 6316
rect 8076 6264 8082 6316
rect 9140 6304 9168 6344
rect 10042 6332 10048 6344
rect 10100 6332 10106 6384
rect 14461 6375 14519 6381
rect 14461 6341 14473 6375
rect 14507 6372 14519 6375
rect 14507 6344 14780 6372
rect 14507 6341 14519 6344
rect 14461 6335 14519 6341
rect 14752 6316 14780 6344
rect 8588 6276 9168 6304
rect 9217 6307 9275 6313
rect 7009 6239 7067 6245
rect 7009 6236 7021 6239
rect 5736 6208 7021 6236
rect 7009 6205 7021 6208
rect 7055 6205 7067 6239
rect 7009 6199 7067 6205
rect 7466 6196 7472 6248
rect 7524 6236 7530 6248
rect 8588 6236 8616 6276
rect 9217 6273 9229 6307
rect 9263 6304 9275 6307
rect 9398 6304 9404 6316
rect 9263 6276 9404 6304
rect 9263 6273 9275 6276
rect 9217 6267 9275 6273
rect 9398 6264 9404 6276
rect 9456 6264 9462 6316
rect 11698 6264 11704 6316
rect 11756 6304 11762 6316
rect 12250 6304 12256 6316
rect 11756 6276 12256 6304
rect 11756 6264 11762 6276
rect 12250 6264 12256 6276
rect 12308 6264 12314 6316
rect 12805 6307 12863 6313
rect 12805 6273 12817 6307
rect 12851 6304 12863 6307
rect 12894 6304 12900 6316
rect 12851 6276 12900 6304
rect 12851 6273 12863 6276
rect 12805 6267 12863 6273
rect 12894 6264 12900 6276
rect 12952 6264 12958 6316
rect 13906 6264 13912 6316
rect 13964 6264 13970 6316
rect 14093 6307 14151 6313
rect 14093 6273 14105 6307
rect 14139 6273 14151 6307
rect 14093 6267 14151 6273
rect 14369 6307 14427 6313
rect 14369 6273 14381 6307
rect 14415 6304 14427 6307
rect 14550 6304 14556 6316
rect 14415 6276 14556 6304
rect 14415 6273 14427 6276
rect 14369 6267 14427 6273
rect 7524 6208 8616 6236
rect 7524 6196 7530 6208
rect 8662 6196 8668 6248
rect 8720 6236 8726 6248
rect 9582 6236 9588 6248
rect 8720 6208 9588 6236
rect 8720 6196 8726 6208
rect 9582 6196 9588 6208
rect 9640 6196 9646 6248
rect 11606 6196 11612 6248
rect 11664 6196 11670 6248
rect 12434 6196 12440 6248
rect 12492 6196 12498 6248
rect 12986 6196 12992 6248
rect 13044 6196 13050 6248
rect 5276 6168 5304 6196
rect 5000 6140 5304 6168
rect 5368 6168 5396 6196
rect 5994 6168 6000 6180
rect 5368 6140 6000 6168
rect 1949 6103 2007 6109
rect 1949 6069 1961 6103
rect 1995 6100 2007 6103
rect 2406 6100 2412 6112
rect 1995 6072 2412 6100
rect 1995 6069 2007 6072
rect 1949 6063 2007 6069
rect 2406 6060 2412 6072
rect 2464 6060 2470 6112
rect 3418 6060 3424 6112
rect 3476 6060 3482 6112
rect 3878 6060 3884 6112
rect 3936 6100 3942 6112
rect 4249 6103 4307 6109
rect 4249 6100 4261 6103
rect 3936 6072 4261 6100
rect 3936 6060 3942 6072
rect 4249 6069 4261 6072
rect 4295 6069 4307 6103
rect 4249 6063 4307 6069
rect 4430 6060 4436 6112
rect 4488 6060 4494 6112
rect 5000 6109 5028 6140
rect 5994 6128 6000 6140
rect 6052 6168 6058 6180
rect 6638 6168 6644 6180
rect 6052 6140 6644 6168
rect 6052 6128 6058 6140
rect 6638 6128 6644 6140
rect 6696 6128 6702 6180
rect 6917 6171 6975 6177
rect 6917 6137 6929 6171
rect 6963 6168 6975 6171
rect 11790 6168 11796 6180
rect 6963 6140 11796 6168
rect 6963 6137 6975 6140
rect 6917 6131 6975 6137
rect 11790 6128 11796 6140
rect 11848 6128 11854 6180
rect 14108 6112 14136 6267
rect 14550 6264 14556 6276
rect 14608 6264 14614 6316
rect 14645 6307 14703 6313
rect 14645 6273 14657 6307
rect 14691 6273 14703 6307
rect 14645 6267 14703 6273
rect 14277 6239 14335 6245
rect 14277 6205 14289 6239
rect 14323 6236 14335 6239
rect 14660 6236 14688 6267
rect 14734 6264 14740 6316
rect 14792 6264 14798 6316
rect 14323 6208 14688 6236
rect 14323 6205 14335 6208
rect 14277 6199 14335 6205
rect 4985 6103 5043 6109
rect 4985 6069 4997 6103
rect 5031 6069 5043 6103
rect 4985 6063 5043 6069
rect 5169 6103 5227 6109
rect 5169 6069 5181 6103
rect 5215 6100 5227 6103
rect 5810 6100 5816 6112
rect 5215 6072 5816 6100
rect 5215 6069 5227 6072
rect 5169 6063 5227 6069
rect 5810 6060 5816 6072
rect 5868 6060 5874 6112
rect 7650 6060 7656 6112
rect 7708 6060 7714 6112
rect 8478 6060 8484 6112
rect 8536 6060 8542 6112
rect 8665 6103 8723 6109
rect 8665 6069 8677 6103
rect 8711 6100 8723 6103
rect 9398 6100 9404 6112
rect 8711 6072 9404 6100
rect 8711 6069 8723 6072
rect 8665 6063 8723 6069
rect 9398 6060 9404 6072
rect 9456 6060 9462 6112
rect 10042 6060 10048 6112
rect 10100 6100 10106 6112
rect 11606 6100 11612 6112
rect 10100 6072 11612 6100
rect 10100 6060 10106 6072
rect 11606 6060 11612 6072
rect 11664 6060 11670 6112
rect 11974 6060 11980 6112
rect 12032 6060 12038 6112
rect 14090 6060 14096 6112
rect 14148 6060 14154 6112
rect 1104 6010 16376 6032
rect 1104 5958 2859 6010
rect 2911 5958 2923 6010
rect 2975 5958 2987 6010
rect 3039 5958 3051 6010
rect 3103 5958 3115 6010
rect 3167 5958 6677 6010
rect 6729 5958 6741 6010
rect 6793 5958 6805 6010
rect 6857 5958 6869 6010
rect 6921 5958 6933 6010
rect 6985 5958 10495 6010
rect 10547 5958 10559 6010
rect 10611 5958 10623 6010
rect 10675 5958 10687 6010
rect 10739 5958 10751 6010
rect 10803 5958 14313 6010
rect 14365 5958 14377 6010
rect 14429 5958 14441 6010
rect 14493 5958 14505 6010
rect 14557 5958 14569 6010
rect 14621 5958 16376 6010
rect 1104 5936 16376 5958
rect 1670 5856 1676 5908
rect 1728 5896 1734 5908
rect 1728 5868 2774 5896
rect 1728 5856 1734 5868
rect 2746 5828 2774 5868
rect 3326 5856 3332 5908
rect 3384 5896 3390 5908
rect 3513 5899 3571 5905
rect 3513 5896 3525 5899
rect 3384 5868 3525 5896
rect 3384 5856 3390 5868
rect 3513 5865 3525 5868
rect 3559 5865 3571 5899
rect 3513 5859 3571 5865
rect 4801 5899 4859 5905
rect 4801 5865 4813 5899
rect 4847 5896 4859 5899
rect 4982 5896 4988 5908
rect 4847 5868 4988 5896
rect 4847 5865 4859 5868
rect 4801 5859 4859 5865
rect 4982 5856 4988 5868
rect 5040 5856 5046 5908
rect 6086 5856 6092 5908
rect 6144 5896 6150 5908
rect 6546 5896 6552 5908
rect 6144 5868 6552 5896
rect 6144 5856 6150 5868
rect 6546 5856 6552 5868
rect 6604 5896 6610 5908
rect 6733 5899 6791 5905
rect 6733 5896 6745 5899
rect 6604 5868 6745 5896
rect 6604 5856 6610 5868
rect 6733 5865 6745 5868
rect 6779 5865 6791 5899
rect 6733 5859 6791 5865
rect 6917 5899 6975 5905
rect 6917 5865 6929 5899
rect 6963 5896 6975 5899
rect 7466 5896 7472 5908
rect 6963 5868 7472 5896
rect 6963 5865 6975 5868
rect 6917 5859 6975 5865
rect 7466 5856 7472 5868
rect 7524 5856 7530 5908
rect 7561 5899 7619 5905
rect 7561 5865 7573 5899
rect 7607 5896 7619 5899
rect 7926 5896 7932 5908
rect 7607 5868 7932 5896
rect 7607 5865 7619 5868
rect 7561 5859 7619 5865
rect 7926 5856 7932 5868
rect 7984 5856 7990 5908
rect 8294 5856 8300 5908
rect 8352 5856 8358 5908
rect 8570 5856 8576 5908
rect 8628 5896 8634 5908
rect 9030 5896 9036 5908
rect 8628 5868 9036 5896
rect 8628 5856 8634 5868
rect 9030 5856 9036 5868
rect 9088 5856 9094 5908
rect 9125 5899 9183 5905
rect 9125 5865 9137 5899
rect 9171 5896 9183 5899
rect 9398 5896 9404 5908
rect 9171 5868 9404 5896
rect 9171 5865 9183 5868
rect 9125 5859 9183 5865
rect 9398 5856 9404 5868
rect 9456 5856 9462 5908
rect 11057 5899 11115 5905
rect 11057 5865 11069 5899
rect 11103 5896 11115 5899
rect 11698 5896 11704 5908
rect 11103 5868 11704 5896
rect 11103 5865 11115 5868
rect 11057 5859 11115 5865
rect 11698 5856 11704 5868
rect 11756 5856 11762 5908
rect 11974 5856 11980 5908
rect 12032 5896 12038 5908
rect 12621 5899 12679 5905
rect 12032 5868 12388 5896
rect 12032 5856 12038 5868
rect 5626 5828 5632 5840
rect 2746 5800 5632 5828
rect 5626 5788 5632 5800
rect 5684 5788 5690 5840
rect 8018 5828 8024 5840
rect 7116 5800 8024 5828
rect 2314 5760 2320 5772
rect 1872 5732 2320 5760
rect 1872 5701 1900 5732
rect 2314 5720 2320 5732
rect 2372 5760 2378 5772
rect 2372 5732 2544 5760
rect 2372 5720 2378 5732
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5661 1639 5695
rect 1857 5695 1915 5701
rect 1857 5692 1869 5695
rect 1581 5655 1639 5661
rect 1688 5664 1869 5692
rect 1596 5556 1624 5655
rect 1688 5636 1716 5664
rect 1857 5661 1869 5664
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 1946 5652 1952 5704
rect 2004 5652 2010 5704
rect 2038 5652 2044 5704
rect 2096 5692 2102 5704
rect 2516 5701 2544 5732
rect 2590 5720 2596 5772
rect 2648 5720 2654 5772
rect 2682 5720 2688 5772
rect 2740 5760 2746 5772
rect 2740 5732 3096 5760
rect 2740 5720 2746 5732
rect 3068 5701 3096 5732
rect 5810 5720 5816 5772
rect 5868 5760 5874 5772
rect 5905 5763 5963 5769
rect 5905 5760 5917 5763
rect 5868 5732 5917 5760
rect 5868 5720 5874 5732
rect 5905 5729 5917 5732
rect 5951 5760 5963 5763
rect 6362 5760 6368 5772
rect 5951 5732 6368 5760
rect 5951 5729 5963 5732
rect 5905 5723 5963 5729
rect 6362 5720 6368 5732
rect 6420 5760 6426 5772
rect 6420 5732 6684 5760
rect 6420 5720 6426 5732
rect 2225 5695 2283 5701
rect 2225 5692 2237 5695
rect 2096 5664 2237 5692
rect 2096 5652 2102 5664
rect 2225 5661 2237 5664
rect 2271 5661 2283 5695
rect 2225 5655 2283 5661
rect 2501 5695 2559 5701
rect 2501 5661 2513 5695
rect 2547 5661 2559 5695
rect 2501 5655 2559 5661
rect 2777 5695 2835 5701
rect 2777 5661 2789 5695
rect 2823 5661 2835 5695
rect 2777 5655 2835 5661
rect 3053 5695 3111 5701
rect 3053 5661 3065 5695
rect 3099 5661 3111 5695
rect 3053 5655 3111 5661
rect 1670 5584 1676 5636
rect 1728 5584 1734 5636
rect 1762 5584 1768 5636
rect 1820 5584 1826 5636
rect 1964 5624 1992 5652
rect 2792 5624 2820 5655
rect 1964 5596 2820 5624
rect 3068 5624 3096 5655
rect 3142 5652 3148 5704
rect 3200 5692 3206 5704
rect 3329 5695 3387 5701
rect 3329 5692 3341 5695
rect 3200 5664 3341 5692
rect 3200 5652 3206 5664
rect 3329 5661 3341 5664
rect 3375 5692 3387 5695
rect 3881 5695 3939 5701
rect 3881 5692 3893 5695
rect 3375 5664 3893 5692
rect 3375 5661 3387 5664
rect 3329 5655 3387 5661
rect 3881 5661 3893 5664
rect 3927 5661 3939 5695
rect 3881 5655 3939 5661
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5692 4123 5695
rect 4154 5692 4160 5704
rect 4111 5664 4160 5692
rect 4111 5661 4123 5664
rect 4065 5655 4123 5661
rect 4154 5652 4160 5664
rect 4212 5652 4218 5704
rect 4522 5652 4528 5704
rect 4580 5692 4586 5704
rect 4580 5664 4752 5692
rect 4580 5652 4586 5664
rect 3973 5627 4031 5633
rect 3068 5596 3128 5624
rect 1854 5556 1860 5568
rect 1596 5528 1860 5556
rect 1854 5516 1860 5528
rect 1912 5516 1918 5568
rect 2130 5516 2136 5568
rect 2188 5516 2194 5568
rect 3100 5556 3128 5596
rect 3973 5593 3985 5627
rect 4019 5624 4031 5627
rect 4430 5624 4436 5636
rect 4019 5596 4436 5624
rect 4019 5593 4031 5596
rect 3973 5587 4031 5593
rect 4430 5584 4436 5596
rect 4488 5624 4494 5636
rect 4617 5627 4675 5633
rect 4617 5624 4629 5627
rect 4488 5596 4629 5624
rect 4488 5584 4494 5596
rect 4617 5593 4629 5596
rect 4663 5593 4675 5627
rect 4724 5624 4752 5664
rect 4798 5652 4804 5704
rect 4856 5652 4862 5704
rect 5994 5652 6000 5704
rect 6052 5652 6058 5704
rect 6086 5652 6092 5704
rect 6144 5652 6150 5704
rect 6178 5652 6184 5704
rect 6236 5652 6242 5704
rect 6196 5624 6224 5652
rect 6549 5627 6607 5633
rect 6549 5624 6561 5627
rect 4724 5596 6224 5624
rect 6288 5596 6561 5624
rect 4617 5587 4675 5593
rect 5994 5556 6000 5568
rect 3100 5528 6000 5556
rect 5994 5516 6000 5528
rect 6052 5556 6058 5568
rect 6288 5556 6316 5596
rect 6549 5593 6561 5596
rect 6595 5593 6607 5627
rect 6656 5624 6684 5732
rect 7116 5701 7144 5800
rect 8018 5788 8024 5800
rect 8076 5788 8082 5840
rect 8312 5828 8340 5856
rect 9309 5831 9367 5837
rect 8312 5800 9260 5828
rect 7193 5763 7251 5769
rect 7193 5729 7205 5763
rect 7239 5760 7251 5763
rect 8386 5760 8392 5772
rect 7239 5732 8392 5760
rect 7239 5729 7251 5732
rect 7193 5723 7251 5729
rect 8386 5720 8392 5732
rect 8444 5760 8450 5772
rect 8444 5732 9076 5760
rect 8444 5720 8450 5732
rect 7101 5695 7159 5701
rect 7101 5661 7113 5695
rect 7147 5661 7159 5695
rect 7101 5655 7159 5661
rect 7285 5695 7343 5701
rect 7285 5661 7297 5695
rect 7331 5692 7343 5695
rect 7377 5695 7435 5701
rect 7377 5692 7389 5695
rect 7331 5664 7389 5692
rect 7331 5661 7343 5664
rect 7285 5655 7343 5661
rect 7377 5661 7389 5664
rect 7423 5692 7435 5695
rect 7650 5692 7656 5704
rect 7423 5664 7656 5692
rect 7423 5661 7435 5664
rect 7377 5655 7435 5661
rect 7650 5652 7656 5664
rect 7708 5652 7714 5704
rect 7926 5652 7932 5704
rect 7984 5692 7990 5704
rect 8021 5695 8079 5701
rect 8021 5692 8033 5695
rect 7984 5664 8033 5692
rect 7984 5652 7990 5664
rect 8021 5661 8033 5664
rect 8067 5661 8079 5695
rect 8021 5655 8079 5661
rect 8478 5652 8484 5704
rect 8536 5692 8542 5704
rect 8536 5664 8984 5692
rect 8536 5652 8542 5664
rect 8956 5633 8984 5664
rect 6749 5627 6807 5633
rect 6749 5624 6761 5627
rect 6656 5596 6761 5624
rect 6549 5587 6607 5593
rect 6749 5593 6761 5596
rect 6795 5593 6807 5627
rect 8941 5627 8999 5633
rect 6749 5587 6807 5593
rect 7484 5596 8892 5624
rect 6052 5528 6316 5556
rect 6365 5559 6423 5565
rect 6052 5516 6058 5528
rect 6365 5525 6377 5559
rect 6411 5556 6423 5559
rect 7484 5556 7512 5596
rect 6411 5528 7512 5556
rect 6411 5525 6423 5528
rect 6365 5519 6423 5525
rect 8202 5516 8208 5568
rect 8260 5516 8266 5568
rect 8294 5516 8300 5568
rect 8352 5556 8358 5568
rect 8570 5556 8576 5568
rect 8352 5528 8576 5556
rect 8352 5516 8358 5528
rect 8570 5516 8576 5528
rect 8628 5516 8634 5568
rect 8864 5556 8892 5596
rect 8941 5593 8953 5627
rect 8987 5593 8999 5627
rect 9048 5624 9076 5732
rect 9141 5627 9199 5633
rect 9141 5624 9153 5627
rect 9048 5596 9153 5624
rect 8941 5587 8999 5593
rect 9141 5593 9153 5596
rect 9187 5593 9199 5627
rect 9232 5624 9260 5800
rect 9309 5797 9321 5831
rect 9355 5797 9367 5831
rect 9309 5791 9367 5797
rect 9953 5831 10011 5837
rect 9953 5797 9965 5831
rect 9999 5797 10011 5831
rect 9953 5791 10011 5797
rect 10597 5831 10655 5837
rect 10597 5797 10609 5831
rect 10643 5828 10655 5831
rect 11514 5828 11520 5840
rect 10643 5800 11520 5828
rect 10643 5797 10655 5800
rect 10597 5791 10655 5797
rect 9324 5760 9352 5791
rect 9493 5763 9551 5769
rect 9493 5760 9505 5763
rect 9324 5732 9505 5760
rect 9493 5729 9505 5732
rect 9539 5729 9551 5763
rect 9493 5723 9551 5729
rect 9582 5652 9588 5704
rect 9640 5652 9646 5704
rect 9968 5692 9996 5791
rect 11514 5788 11520 5800
rect 11572 5788 11578 5840
rect 11606 5788 11612 5840
rect 11664 5828 11670 5840
rect 12115 5831 12173 5837
rect 12115 5828 12127 5831
rect 11664 5800 12127 5828
rect 11664 5788 11670 5800
rect 12115 5797 12127 5800
rect 12161 5797 12173 5831
rect 12115 5791 12173 5797
rect 12360 5769 12388 5868
rect 12621 5865 12633 5899
rect 12667 5896 12679 5899
rect 12986 5896 12992 5908
rect 12667 5868 12992 5896
rect 12667 5865 12679 5868
rect 12621 5859 12679 5865
rect 12986 5856 12992 5868
rect 13044 5856 13050 5908
rect 14642 5856 14648 5908
rect 14700 5856 14706 5908
rect 10689 5763 10747 5769
rect 10689 5760 10701 5763
rect 10428 5732 10701 5760
rect 10428 5701 10456 5732
rect 10689 5729 10701 5732
rect 10735 5729 10747 5763
rect 12345 5763 12403 5769
rect 12345 5760 12357 5763
rect 10689 5723 10747 5729
rect 11440 5732 12357 5760
rect 11440 5701 11468 5732
rect 12345 5729 12357 5732
rect 12391 5729 12403 5763
rect 12345 5723 12403 5729
rect 13817 5763 13875 5769
rect 13817 5729 13829 5763
rect 13863 5760 13875 5763
rect 14090 5760 14096 5772
rect 13863 5732 14096 5760
rect 13863 5729 13875 5732
rect 13817 5723 13875 5729
rect 14090 5720 14096 5732
rect 14148 5760 14154 5772
rect 14185 5763 14243 5769
rect 14185 5760 14197 5763
rect 14148 5732 14197 5760
rect 14148 5720 14154 5732
rect 14185 5729 14197 5732
rect 14231 5729 14243 5763
rect 14660 5760 14688 5856
rect 14829 5763 14887 5769
rect 14829 5760 14841 5763
rect 14660 5732 14841 5760
rect 14185 5723 14243 5729
rect 14829 5729 14841 5732
rect 14875 5729 14887 5763
rect 14829 5723 14887 5729
rect 15289 5763 15347 5769
rect 15289 5729 15301 5763
rect 15335 5760 15347 5763
rect 15335 5732 15700 5760
rect 15335 5729 15347 5732
rect 15289 5723 15347 5729
rect 10413 5695 10471 5701
rect 10413 5692 10425 5695
rect 9968 5664 10425 5692
rect 10413 5661 10425 5664
rect 10459 5661 10471 5695
rect 10413 5655 10471 5661
rect 10597 5695 10655 5701
rect 10597 5661 10609 5695
rect 10643 5692 10655 5695
rect 10873 5695 10931 5701
rect 10873 5692 10885 5695
rect 10643 5664 10885 5692
rect 10643 5661 10655 5664
rect 10597 5655 10655 5661
rect 10873 5661 10885 5664
rect 10919 5661 10931 5695
rect 10873 5655 10931 5661
rect 11425 5695 11483 5701
rect 11425 5661 11437 5695
rect 11471 5661 11483 5695
rect 11425 5655 11483 5661
rect 11517 5695 11575 5701
rect 11517 5661 11529 5695
rect 11563 5661 11575 5695
rect 11517 5655 11575 5661
rect 11701 5695 11759 5701
rect 11701 5661 11713 5695
rect 11747 5692 11759 5695
rect 11790 5692 11796 5704
rect 11747 5664 11796 5692
rect 11747 5661 11759 5664
rect 11701 5655 11759 5661
rect 10612 5624 10640 5655
rect 9232 5596 10640 5624
rect 11532 5624 11560 5655
rect 11790 5652 11796 5664
rect 11848 5692 11854 5704
rect 12207 5695 12265 5701
rect 12207 5692 12219 5695
rect 11848 5664 12219 5692
rect 11848 5652 11854 5664
rect 12207 5661 12219 5664
rect 12253 5661 12265 5695
rect 12207 5655 12265 5661
rect 12894 5652 12900 5704
rect 12952 5692 12958 5704
rect 13081 5695 13139 5701
rect 13081 5692 13093 5695
rect 12952 5664 13093 5692
rect 12952 5652 12958 5664
rect 13081 5661 13093 5664
rect 13127 5661 13139 5695
rect 13081 5655 13139 5661
rect 13354 5652 13360 5704
rect 13412 5652 13418 5704
rect 13906 5652 13912 5704
rect 13964 5692 13970 5704
rect 14277 5695 14335 5701
rect 14277 5692 14289 5695
rect 13964 5664 14289 5692
rect 13964 5652 13970 5664
rect 14277 5661 14289 5664
rect 14323 5661 14335 5695
rect 14277 5655 14335 5661
rect 14734 5652 14740 5704
rect 14792 5692 14798 5704
rect 15672 5701 15700 5732
rect 14921 5695 14979 5701
rect 14921 5692 14933 5695
rect 14792 5664 14933 5692
rect 14792 5652 14798 5664
rect 14921 5661 14933 5664
rect 14967 5661 14979 5695
rect 14921 5655 14979 5661
rect 15657 5695 15715 5701
rect 15657 5661 15669 5695
rect 15703 5661 15715 5695
rect 15657 5655 15715 5661
rect 11977 5627 12035 5633
rect 11977 5624 11989 5627
rect 11532 5596 11989 5624
rect 9141 5587 9199 5593
rect 11624 5568 11652 5596
rect 11977 5593 11989 5596
rect 12023 5593 12035 5627
rect 11977 5587 12035 5593
rect 9674 5556 9680 5568
rect 8864 5528 9680 5556
rect 9674 5516 9680 5528
rect 9732 5516 9738 5568
rect 11606 5516 11612 5568
rect 11664 5516 11670 5568
rect 11885 5559 11943 5565
rect 11885 5525 11897 5559
rect 11931 5556 11943 5559
rect 12434 5556 12440 5568
rect 11931 5528 12440 5556
rect 11931 5525 11943 5528
rect 11885 5519 11943 5525
rect 12434 5516 12440 5528
rect 12492 5556 12498 5568
rect 13170 5556 13176 5568
rect 12492 5528 13176 5556
rect 12492 5516 12498 5528
rect 13170 5516 13176 5528
rect 13228 5516 13234 5568
rect 15933 5559 15991 5565
rect 15933 5525 15945 5559
rect 15979 5556 15991 5559
rect 16022 5556 16028 5568
rect 15979 5528 16028 5556
rect 15979 5525 15991 5528
rect 15933 5519 15991 5525
rect 16022 5516 16028 5528
rect 16080 5516 16086 5568
rect 1104 5466 16376 5488
rect 1104 5414 3519 5466
rect 3571 5414 3583 5466
rect 3635 5414 3647 5466
rect 3699 5414 3711 5466
rect 3763 5414 3775 5466
rect 3827 5414 7337 5466
rect 7389 5414 7401 5466
rect 7453 5414 7465 5466
rect 7517 5414 7529 5466
rect 7581 5414 7593 5466
rect 7645 5414 11155 5466
rect 11207 5414 11219 5466
rect 11271 5414 11283 5466
rect 11335 5414 11347 5466
rect 11399 5414 11411 5466
rect 11463 5414 14973 5466
rect 15025 5414 15037 5466
rect 15089 5414 15101 5466
rect 15153 5414 15165 5466
rect 15217 5414 15229 5466
rect 15281 5414 16376 5466
rect 1104 5392 16376 5414
rect 4338 5312 4344 5364
rect 4396 5312 4402 5364
rect 4522 5312 4528 5364
rect 4580 5312 4586 5364
rect 8386 5312 8392 5364
rect 8444 5312 8450 5364
rect 8478 5312 8484 5364
rect 8536 5352 8542 5364
rect 8536 5324 9260 5352
rect 8536 5312 8542 5324
rect 2409 5287 2467 5293
rect 2409 5253 2421 5287
rect 2455 5284 2467 5287
rect 2498 5284 2504 5296
rect 2455 5256 2504 5284
rect 2455 5253 2467 5256
rect 2409 5247 2467 5253
rect 2498 5244 2504 5256
rect 2556 5244 2562 5296
rect 2685 5287 2743 5293
rect 2685 5253 2697 5287
rect 2731 5284 2743 5287
rect 2774 5284 2780 5296
rect 2731 5256 2780 5284
rect 2731 5253 2743 5256
rect 2685 5247 2743 5253
rect 2774 5244 2780 5256
rect 2832 5244 2838 5296
rect 2869 5287 2927 5293
rect 2869 5253 2881 5287
rect 2915 5284 2927 5287
rect 3142 5284 3148 5296
rect 2915 5256 3148 5284
rect 2915 5253 2927 5256
rect 2869 5247 2927 5253
rect 3142 5244 3148 5256
rect 3200 5244 3206 5296
rect 1670 5176 1676 5228
rect 1728 5216 1734 5228
rect 1857 5219 1915 5225
rect 1857 5216 1869 5219
rect 1728 5188 1869 5216
rect 1728 5176 1734 5188
rect 1857 5185 1869 5188
rect 1903 5185 1915 5219
rect 1857 5179 1915 5185
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5185 4215 5219
rect 4157 5179 4215 5185
rect 2590 5108 2596 5160
rect 2648 5148 2654 5160
rect 3510 5148 3516 5160
rect 2648 5120 3516 5148
rect 2648 5108 2654 5120
rect 3510 5108 3516 5120
rect 3568 5148 3574 5160
rect 3789 5151 3847 5157
rect 3789 5148 3801 5151
rect 3568 5120 3801 5148
rect 3568 5108 3574 5120
rect 3789 5117 3801 5120
rect 3835 5117 3847 5151
rect 3789 5111 3847 5117
rect 4172 5024 4200 5179
rect 4246 5176 4252 5228
rect 4304 5216 4310 5228
rect 4356 5216 4384 5312
rect 4540 5284 4568 5312
rect 4448 5256 4568 5284
rect 4448 5225 4476 5256
rect 7834 5244 7840 5296
rect 7892 5244 7898 5296
rect 7926 5244 7932 5296
rect 7984 5244 7990 5296
rect 8404 5284 8432 5312
rect 8404 5256 9168 5284
rect 5080 5228 5132 5234
rect 4304 5188 4384 5216
rect 4433 5219 4491 5225
rect 4304 5176 4310 5188
rect 4433 5185 4445 5219
rect 4479 5185 4491 5219
rect 4433 5179 4491 5185
rect 6362 5176 6368 5228
rect 6420 5176 6426 5228
rect 6641 5219 6699 5225
rect 6641 5185 6653 5219
rect 6687 5216 6699 5219
rect 7469 5219 7527 5225
rect 7469 5216 7481 5219
rect 6687 5188 7481 5216
rect 6687 5185 6699 5188
rect 6641 5179 6699 5185
rect 7469 5185 7481 5188
rect 7515 5185 7527 5219
rect 7469 5179 7527 5185
rect 7653 5219 7711 5225
rect 7653 5185 7665 5219
rect 7699 5185 7711 5219
rect 7653 5179 7711 5185
rect 8021 5219 8079 5225
rect 8021 5185 8033 5219
rect 8067 5216 8079 5219
rect 8294 5216 8300 5228
rect 8067 5188 8300 5216
rect 8067 5185 8079 5188
rect 8021 5179 8079 5185
rect 5080 5170 5132 5176
rect 5350 5108 5356 5160
rect 5408 5108 5414 5160
rect 7668 5148 7696 5179
rect 8294 5176 8300 5188
rect 8352 5176 8358 5228
rect 8404 5216 8432 5256
rect 8481 5219 8539 5225
rect 8481 5216 8493 5219
rect 8404 5188 8493 5216
rect 8481 5185 8493 5188
rect 8527 5185 8539 5219
rect 8481 5179 8539 5185
rect 8573 5219 8631 5225
rect 8573 5185 8585 5219
rect 8619 5216 8631 5219
rect 8662 5216 8668 5228
rect 8619 5188 8668 5216
rect 8619 5185 8631 5188
rect 8573 5179 8631 5185
rect 8662 5176 8668 5188
rect 8720 5176 8726 5228
rect 9140 5225 9168 5256
rect 9232 5225 9260 5324
rect 9674 5312 9680 5364
rect 9732 5312 9738 5364
rect 13265 5355 13323 5361
rect 13265 5321 13277 5355
rect 13311 5352 13323 5355
rect 13354 5352 13360 5364
rect 13311 5324 13360 5352
rect 13311 5321 13323 5324
rect 13265 5315 13323 5321
rect 13354 5312 13360 5324
rect 13412 5312 13418 5364
rect 8757 5219 8815 5225
rect 8757 5185 8769 5219
rect 8803 5216 8815 5219
rect 9125 5219 9183 5225
rect 8803 5188 9076 5216
rect 8803 5185 8815 5188
rect 8757 5179 8815 5185
rect 8386 5148 8392 5160
rect 7668 5120 8392 5148
rect 8386 5108 8392 5120
rect 8444 5108 8450 5160
rect 8849 5151 8907 5157
rect 8849 5117 8861 5151
rect 8895 5117 8907 5151
rect 8849 5111 8907 5117
rect 8205 5083 8263 5089
rect 8205 5049 8217 5083
rect 8251 5080 8263 5083
rect 8864 5080 8892 5111
rect 9048 5089 9076 5188
rect 9125 5185 9137 5219
rect 9171 5185 9183 5219
rect 9125 5179 9183 5185
rect 9217 5219 9275 5225
rect 9217 5185 9229 5219
rect 9263 5185 9275 5219
rect 9217 5179 9275 5185
rect 9394 5219 9452 5225
rect 9394 5185 9406 5219
rect 9440 5185 9452 5219
rect 9692 5216 9720 5312
rect 11514 5244 11520 5296
rect 11572 5244 11578 5296
rect 11698 5244 11704 5296
rect 11756 5244 11762 5296
rect 9953 5219 10011 5225
rect 9953 5216 9965 5219
rect 9692 5188 9965 5216
rect 9394 5179 9452 5185
rect 9953 5185 9965 5188
rect 9999 5185 10011 5219
rect 9953 5179 10011 5185
rect 10781 5219 10839 5225
rect 10781 5185 10793 5219
rect 10827 5216 10839 5219
rect 12805 5219 12863 5225
rect 10827 5188 11284 5216
rect 10827 5185 10839 5188
rect 10781 5179 10839 5185
rect 9416 5092 9444 5179
rect 8251 5052 8892 5080
rect 9033 5083 9091 5089
rect 8251 5049 8263 5052
rect 8205 5043 8263 5049
rect 9033 5049 9045 5083
rect 9079 5080 9091 5083
rect 9309 5083 9367 5089
rect 9309 5080 9321 5083
rect 9079 5052 9321 5080
rect 9079 5049 9091 5052
rect 9033 5043 9091 5049
rect 9309 5049 9321 5052
rect 9355 5049 9367 5083
rect 9309 5043 9367 5049
rect 9398 5040 9404 5092
rect 9456 5040 9462 5092
rect 11256 5024 11284 5188
rect 12805 5185 12817 5219
rect 12851 5216 12863 5219
rect 12986 5216 12992 5228
rect 12851 5188 12992 5216
rect 12851 5185 12863 5188
rect 12805 5179 12863 5185
rect 12986 5176 12992 5188
rect 13044 5176 13050 5228
rect 13170 5176 13176 5228
rect 13228 5176 13234 5228
rect 3970 4972 3976 5024
rect 4028 4972 4034 5024
rect 4154 4972 4160 5024
rect 4212 4972 4218 5024
rect 6086 4972 6092 5024
rect 6144 5012 6150 5024
rect 7285 5015 7343 5021
rect 7285 5012 7297 5015
rect 6144 4984 7297 5012
rect 6144 4972 6150 4984
rect 7285 4981 7297 4984
rect 7331 4981 7343 5015
rect 7285 4975 7343 4981
rect 8754 4972 8760 5024
rect 8812 4972 8818 5024
rect 8938 4972 8944 5024
rect 8996 4972 9002 5024
rect 10042 4972 10048 5024
rect 10100 4972 10106 5024
rect 10410 4972 10416 5024
rect 10468 4972 10474 5024
rect 10597 5015 10655 5021
rect 10597 4981 10609 5015
rect 10643 5012 10655 5015
rect 10870 5012 10876 5024
rect 10643 4984 10876 5012
rect 10643 4981 10655 4984
rect 10597 4975 10655 4981
rect 10870 4972 10876 4984
rect 10928 4972 10934 5024
rect 11238 4972 11244 5024
rect 11296 4972 11302 5024
rect 11882 4972 11888 5024
rect 11940 4972 11946 5024
rect 1104 4922 16376 4944
rect 1104 4870 2859 4922
rect 2911 4870 2923 4922
rect 2975 4870 2987 4922
rect 3039 4870 3051 4922
rect 3103 4870 3115 4922
rect 3167 4870 6677 4922
rect 6729 4870 6741 4922
rect 6793 4870 6805 4922
rect 6857 4870 6869 4922
rect 6921 4870 6933 4922
rect 6985 4870 10495 4922
rect 10547 4870 10559 4922
rect 10611 4870 10623 4922
rect 10675 4870 10687 4922
rect 10739 4870 10751 4922
rect 10803 4870 14313 4922
rect 14365 4870 14377 4922
rect 14429 4870 14441 4922
rect 14493 4870 14505 4922
rect 14557 4870 14569 4922
rect 14621 4870 16376 4922
rect 1104 4848 16376 4870
rect 2961 4811 3019 4817
rect 2961 4808 2973 4811
rect 2240 4780 2973 4808
rect 1762 4632 1768 4684
rect 1820 4632 1826 4684
rect 934 4564 940 4616
rect 992 4604 998 4616
rect 1489 4607 1547 4613
rect 1489 4604 1501 4607
rect 992 4576 1501 4604
rect 992 4564 998 4576
rect 1489 4573 1501 4576
rect 1535 4573 1547 4607
rect 1489 4567 1547 4573
rect 2130 4564 2136 4616
rect 2188 4604 2194 4616
rect 2240 4613 2268 4780
rect 2961 4777 2973 4780
rect 3007 4808 3019 4811
rect 3007 4780 3464 4808
rect 3007 4777 3019 4780
rect 2961 4771 3019 4777
rect 2685 4675 2743 4681
rect 2685 4641 2697 4675
rect 2731 4672 2743 4675
rect 2774 4672 2780 4684
rect 2731 4644 2780 4672
rect 2731 4641 2743 4644
rect 2685 4635 2743 4641
rect 2774 4632 2780 4644
rect 2832 4632 2838 4684
rect 2225 4607 2283 4613
rect 2225 4604 2237 4607
rect 2188 4576 2237 4604
rect 2188 4564 2194 4576
rect 2225 4573 2237 4576
rect 2271 4573 2283 4607
rect 2225 4567 2283 4573
rect 2406 4564 2412 4616
rect 2464 4604 2470 4616
rect 3436 4613 3464 4780
rect 3510 4768 3516 4820
rect 3568 4768 3574 4820
rect 3970 4768 3976 4820
rect 4028 4768 4034 4820
rect 5997 4811 6055 4817
rect 5997 4777 6009 4811
rect 6043 4808 6055 4811
rect 7006 4808 7012 4820
rect 6043 4780 7012 4808
rect 6043 4777 6055 4780
rect 5997 4771 6055 4777
rect 3528 4613 3556 4768
rect 3988 4672 4016 4768
rect 6086 4700 6092 4752
rect 6144 4700 6150 4752
rect 5813 4675 5871 4681
rect 5813 4672 5825 4675
rect 3988 4644 5825 4672
rect 5813 4641 5825 4644
rect 5859 4641 5871 4675
rect 5813 4635 5871 4641
rect 2501 4607 2559 4613
rect 2501 4604 2513 4607
rect 2464 4576 2513 4604
rect 2464 4564 2470 4576
rect 2501 4573 2513 4576
rect 2547 4604 2559 4607
rect 3237 4607 3295 4613
rect 3237 4604 3249 4607
rect 2547 4576 3249 4604
rect 2547 4573 2559 4576
rect 2501 4567 2559 4573
rect 2317 4539 2375 4545
rect 2317 4505 2329 4539
rect 2363 4536 2375 4539
rect 2590 4536 2596 4548
rect 2363 4508 2596 4536
rect 2363 4505 2375 4508
rect 2317 4499 2375 4505
rect 2590 4496 2596 4508
rect 2648 4536 2654 4548
rect 2976 4545 3004 4576
rect 3237 4573 3249 4576
rect 3283 4573 3295 4607
rect 3237 4567 3295 4573
rect 3421 4607 3479 4613
rect 3421 4573 3433 4607
rect 3467 4573 3479 4607
rect 3421 4567 3479 4573
rect 3513 4607 3571 4613
rect 3513 4573 3525 4607
rect 3559 4573 3571 4607
rect 3513 4567 3571 4573
rect 4154 4564 4160 4616
rect 4212 4564 4218 4616
rect 2777 4539 2835 4545
rect 2777 4536 2789 4539
rect 2648 4508 2789 4536
rect 2648 4496 2654 4508
rect 2777 4505 2789 4508
rect 2823 4505 2835 4539
rect 2976 4539 3035 4545
rect 2976 4508 2989 4539
rect 2777 4499 2835 4505
rect 2977 4505 2989 4508
rect 3023 4505 3035 4539
rect 4172 4536 4200 4564
rect 2977 4499 3035 4505
rect 3160 4508 4200 4536
rect 5828 4536 5856 4635
rect 6104 4613 6132 4700
rect 6196 4613 6224 4780
rect 7006 4768 7012 4780
rect 7064 4768 7070 4820
rect 10410 4768 10416 4820
rect 10468 4768 10474 4820
rect 10870 4768 10876 4820
rect 10928 4768 10934 4820
rect 11425 4811 11483 4817
rect 11425 4777 11437 4811
rect 11471 4808 11483 4811
rect 11606 4808 11612 4820
rect 11471 4780 11612 4808
rect 11471 4777 11483 4780
rect 11425 4771 11483 4777
rect 11606 4768 11612 4780
rect 11664 4768 11670 4820
rect 6273 4743 6331 4749
rect 6273 4709 6285 4743
rect 6319 4740 6331 4743
rect 6362 4740 6368 4752
rect 6319 4712 6368 4740
rect 6319 4709 6331 4712
rect 6273 4703 6331 4709
rect 6362 4700 6368 4712
rect 6420 4700 6426 4752
rect 7469 4675 7527 4681
rect 7469 4641 7481 4675
rect 7515 4672 7527 4675
rect 7650 4672 7656 4684
rect 7515 4644 7656 4672
rect 7515 4641 7527 4644
rect 7469 4635 7527 4641
rect 7650 4632 7656 4644
rect 7708 4672 7714 4684
rect 10428 4681 10456 4768
rect 10888 4740 10916 4768
rect 10520 4712 10916 4740
rect 8297 4675 8355 4681
rect 8297 4672 8309 4675
rect 7708 4644 8309 4672
rect 7708 4632 7714 4644
rect 8297 4641 8309 4644
rect 8343 4641 8355 4675
rect 8297 4635 8355 4641
rect 10413 4675 10471 4681
rect 10413 4641 10425 4675
rect 10459 4641 10471 4675
rect 10413 4635 10471 4641
rect 6089 4607 6147 4613
rect 6089 4573 6101 4607
rect 6135 4573 6147 4607
rect 6089 4567 6147 4573
rect 6181 4607 6239 4613
rect 6181 4573 6193 4607
rect 6227 4573 6239 4607
rect 6181 4567 6239 4573
rect 6457 4607 6515 4613
rect 6457 4573 6469 4607
rect 6503 4573 6515 4607
rect 6457 4567 6515 4573
rect 6472 4536 6500 4567
rect 7098 4564 7104 4616
rect 7156 4604 7162 4616
rect 7377 4607 7435 4613
rect 7377 4604 7389 4607
rect 7156 4576 7389 4604
rect 7156 4564 7162 4576
rect 7377 4573 7389 4576
rect 7423 4573 7435 4607
rect 7377 4567 7435 4573
rect 7558 4564 7564 4616
rect 7616 4604 7622 4616
rect 7745 4607 7803 4613
rect 7745 4604 7757 4607
rect 7616 4576 7757 4604
rect 7616 4564 7622 4576
rect 7745 4573 7757 4576
rect 7791 4573 7803 4607
rect 7745 4567 7803 4573
rect 7837 4607 7895 4613
rect 7837 4573 7849 4607
rect 7883 4573 7895 4607
rect 7837 4567 7895 4573
rect 5828 4508 6500 4536
rect 6917 4539 6975 4545
rect 3160 4477 3188 4508
rect 6917 4505 6929 4539
rect 6963 4536 6975 4539
rect 7009 4539 7067 4545
rect 7009 4536 7021 4539
rect 6963 4508 7021 4536
rect 6963 4505 6975 4508
rect 6917 4499 6975 4505
rect 7009 4505 7021 4508
rect 7055 4536 7067 4539
rect 7852 4536 7880 4567
rect 7055 4508 7880 4536
rect 10428 4536 10456 4635
rect 10520 4613 10548 4712
rect 11238 4700 11244 4752
rect 11296 4700 11302 4752
rect 10873 4675 10931 4681
rect 10873 4641 10885 4675
rect 10919 4672 10931 4675
rect 11054 4672 11060 4684
rect 10919 4644 11060 4672
rect 10919 4641 10931 4644
rect 10873 4635 10931 4641
rect 11054 4632 11060 4644
rect 11112 4632 11118 4684
rect 10505 4607 10563 4613
rect 10505 4573 10517 4607
rect 10551 4573 10563 4607
rect 10505 4567 10563 4573
rect 10965 4539 11023 4545
rect 10965 4536 10977 4539
rect 10428 4508 10977 4536
rect 7055 4505 7067 4508
rect 7009 4499 7067 4505
rect 10965 4505 10977 4508
rect 11011 4505 11023 4539
rect 10965 4499 11023 4505
rect 3145 4471 3203 4477
rect 3145 4437 3157 4471
rect 3191 4437 3203 4471
rect 3145 4431 3203 4437
rect 3326 4428 3332 4480
rect 3384 4428 3390 4480
rect 4338 4428 4344 4480
rect 4396 4428 4402 4480
rect 5813 4471 5871 4477
rect 5813 4437 5825 4471
rect 5859 4468 5871 4471
rect 7558 4468 7564 4480
rect 5859 4440 7564 4468
rect 5859 4437 5871 4440
rect 5813 4431 5871 4437
rect 7558 4428 7564 4440
rect 7616 4428 7622 4480
rect 7653 4471 7711 4477
rect 7653 4437 7665 4471
rect 7699 4468 7711 4471
rect 11256 4468 11284 4700
rect 7699 4440 11284 4468
rect 7699 4437 7711 4440
rect 7653 4431 7711 4437
rect 1104 4378 16376 4400
rect 1104 4326 3519 4378
rect 3571 4326 3583 4378
rect 3635 4326 3647 4378
rect 3699 4326 3711 4378
rect 3763 4326 3775 4378
rect 3827 4326 7337 4378
rect 7389 4326 7401 4378
rect 7453 4326 7465 4378
rect 7517 4326 7529 4378
rect 7581 4326 7593 4378
rect 7645 4326 11155 4378
rect 11207 4326 11219 4378
rect 11271 4326 11283 4378
rect 11335 4326 11347 4378
rect 11399 4326 11411 4378
rect 11463 4326 14973 4378
rect 15025 4326 15037 4378
rect 15089 4326 15101 4378
rect 15153 4326 15165 4378
rect 15217 4326 15229 4378
rect 15281 4326 16376 4378
rect 1104 4304 16376 4326
rect 1854 4224 1860 4276
rect 1912 4264 1918 4276
rect 2133 4267 2191 4273
rect 2133 4264 2145 4267
rect 1912 4236 2145 4264
rect 1912 4224 1918 4236
rect 2133 4233 2145 4236
rect 2179 4233 2191 4267
rect 3605 4267 3663 4273
rect 3605 4264 3617 4267
rect 2133 4227 2191 4233
rect 2792 4236 3617 4264
rect 2792 4208 2820 4236
rect 3605 4233 3617 4236
rect 3651 4233 3663 4267
rect 3605 4227 3663 4233
rect 3878 4224 3884 4276
rect 3936 4224 3942 4276
rect 4890 4224 4896 4276
rect 4948 4224 4954 4276
rect 1026 4156 1032 4208
rect 1084 4196 1090 4208
rect 2041 4199 2099 4205
rect 2041 4196 2053 4199
rect 1084 4168 2053 4196
rect 1084 4156 1090 4168
rect 2041 4165 2053 4168
rect 2087 4165 2099 4199
rect 2041 4159 2099 4165
rect 2774 4156 2780 4208
rect 2832 4156 2838 4208
rect 2869 4199 2927 4205
rect 2869 4165 2881 4199
rect 2915 4196 2927 4199
rect 3237 4199 3295 4205
rect 2915 4168 3188 4196
rect 2915 4165 2927 4168
rect 2869 4159 2927 4165
rect 1394 4088 1400 4140
rect 1452 4088 1458 4140
rect 1670 4088 1676 4140
rect 1728 4088 1734 4140
rect 2593 4131 2651 4137
rect 2593 4097 2605 4131
rect 2639 4128 2651 4131
rect 2961 4131 3019 4137
rect 2639 4100 2728 4128
rect 2639 4097 2651 4100
rect 2593 4091 2651 4097
rect 2700 3992 2728 4100
rect 2961 4097 2973 4131
rect 3007 4097 3019 4131
rect 3160 4128 3188 4168
rect 3237 4165 3249 4199
rect 3283 4196 3295 4199
rect 3326 4196 3332 4208
rect 3283 4168 3332 4196
rect 3283 4165 3295 4168
rect 3237 4159 3295 4165
rect 3326 4156 3332 4168
rect 3384 4156 3390 4208
rect 3421 4199 3479 4205
rect 3421 4165 3433 4199
rect 3467 4196 3479 4199
rect 3896 4196 3924 4224
rect 4908 4196 4936 4224
rect 3467 4168 3924 4196
rect 3988 4168 4936 4196
rect 12360 4168 12664 4196
rect 3467 4165 3479 4168
rect 3421 4159 3479 4165
rect 3436 4128 3464 4159
rect 3160 4100 3464 4128
rect 3513 4131 3571 4137
rect 2961 4091 3019 4097
rect 3513 4097 3525 4131
rect 3559 4128 3571 4131
rect 3988 4128 4016 4168
rect 3559 4100 4016 4128
rect 3559 4097 3571 4100
rect 3513 4091 3571 4097
rect 2976 4060 3004 4091
rect 3528 4060 3556 4091
rect 4062 4088 4068 4140
rect 4120 4088 4126 4140
rect 4157 4131 4215 4137
rect 4157 4097 4169 4131
rect 4203 4128 4215 4131
rect 4338 4128 4344 4140
rect 4203 4100 4344 4128
rect 4203 4097 4215 4100
rect 4157 4091 4215 4097
rect 4338 4088 4344 4100
rect 4396 4088 4402 4140
rect 7006 4088 7012 4140
rect 7064 4128 7070 4140
rect 7377 4131 7435 4137
rect 7377 4128 7389 4131
rect 7064 4100 7389 4128
rect 7064 4088 7070 4100
rect 7377 4097 7389 4100
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 8757 4131 8815 4137
rect 8757 4097 8769 4131
rect 8803 4128 8815 4131
rect 8938 4128 8944 4140
rect 8803 4100 8944 4128
rect 8803 4097 8815 4100
rect 8757 4091 8815 4097
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 9217 4131 9275 4137
rect 9217 4097 9229 4131
rect 9263 4097 9275 4131
rect 9217 4091 9275 4097
rect 2976 4032 3556 4060
rect 3234 3992 3240 4004
rect 2700 3964 3240 3992
rect 3234 3952 3240 3964
rect 3292 3952 3298 4004
rect 4080 3992 4108 4088
rect 4246 4020 4252 4072
rect 4304 4020 4310 4072
rect 7469 4063 7527 4069
rect 7469 4029 7481 4063
rect 7515 4060 7527 4063
rect 7650 4060 7656 4072
rect 7515 4032 7656 4060
rect 7515 4029 7527 4032
rect 7469 4023 7527 4029
rect 7650 4020 7656 4032
rect 7708 4020 7714 4072
rect 7745 4063 7803 4069
rect 7745 4029 7757 4063
rect 7791 4060 7803 4063
rect 8665 4063 8723 4069
rect 8665 4060 8677 4063
rect 7791 4032 8677 4060
rect 7791 4029 7803 4032
rect 7745 4023 7803 4029
rect 8665 4029 8677 4032
rect 8711 4060 8723 4063
rect 9232 4060 9260 4091
rect 11054 4088 11060 4140
rect 11112 4128 11118 4140
rect 11517 4131 11575 4137
rect 11517 4128 11529 4131
rect 11112 4100 11529 4128
rect 11112 4088 11118 4100
rect 11517 4097 11529 4100
rect 11563 4097 11575 4131
rect 11517 4091 11575 4097
rect 11701 4131 11759 4137
rect 11701 4097 11713 4131
rect 11747 4128 11759 4131
rect 11882 4128 11888 4140
rect 11747 4100 11888 4128
rect 11747 4097 11759 4100
rect 11701 4091 11759 4097
rect 8711 4032 9260 4060
rect 11532 4060 11560 4091
rect 11882 4088 11888 4100
rect 11940 4128 11946 4140
rect 11977 4131 12035 4137
rect 11977 4128 11989 4131
rect 11940 4100 11989 4128
rect 11940 4088 11946 4100
rect 11977 4097 11989 4100
rect 12023 4097 12035 4131
rect 11977 4091 12035 4097
rect 12069 4063 12127 4069
rect 12069 4060 12081 4063
rect 11532 4032 12081 4060
rect 8711 4029 8723 4032
rect 8665 4023 8723 4029
rect 12069 4029 12081 4032
rect 12115 4029 12127 4063
rect 12069 4023 12127 4029
rect 8294 3992 8300 4004
rect 4080 3964 8300 3992
rect 8294 3952 8300 3964
rect 8352 3952 8358 4004
rect 11517 3995 11575 4001
rect 8956 3964 9260 3992
rect 8956 3936 8984 3964
rect 3145 3927 3203 3933
rect 3145 3893 3157 3927
rect 3191 3924 3203 3927
rect 3326 3924 3332 3936
rect 3191 3896 3332 3924
rect 3191 3893 3203 3896
rect 3145 3887 3203 3893
rect 3326 3884 3332 3896
rect 3384 3884 3390 3936
rect 3789 3927 3847 3933
rect 3789 3893 3801 3927
rect 3835 3924 3847 3927
rect 3970 3924 3976 3936
rect 3835 3896 3976 3924
rect 3835 3893 3847 3896
rect 3789 3887 3847 3893
rect 3970 3884 3976 3896
rect 4028 3884 4034 3936
rect 4430 3884 4436 3936
rect 4488 3884 4494 3936
rect 7190 3884 7196 3936
rect 7248 3924 7254 3936
rect 8110 3924 8116 3936
rect 7248 3896 8116 3924
rect 7248 3884 7254 3896
rect 8110 3884 8116 3896
rect 8168 3884 8174 3936
rect 8938 3884 8944 3936
rect 8996 3884 9002 3936
rect 9122 3884 9128 3936
rect 9180 3884 9186 3936
rect 9232 3924 9260 3964
rect 11517 3961 11529 3995
rect 11563 3992 11575 3995
rect 12360 3992 12388 4168
rect 12437 4131 12495 4137
rect 12437 4097 12449 4131
rect 12483 4097 12495 4131
rect 12437 4091 12495 4097
rect 12529 4131 12587 4137
rect 12529 4097 12541 4131
rect 12575 4097 12587 4131
rect 12636 4128 12664 4168
rect 12713 4131 12771 4137
rect 12713 4128 12725 4131
rect 12636 4100 12725 4128
rect 12529 4091 12587 4097
rect 12713 4097 12725 4100
rect 12759 4097 12771 4131
rect 12713 4091 12771 4097
rect 11563 3964 12388 3992
rect 11563 3961 11575 3964
rect 11517 3955 11575 3961
rect 9309 3927 9367 3933
rect 9309 3924 9321 3927
rect 9232 3896 9321 3924
rect 9309 3893 9321 3896
rect 9355 3893 9367 3927
rect 9309 3887 9367 3893
rect 9674 3884 9680 3936
rect 9732 3884 9738 3936
rect 12345 3927 12403 3933
rect 12345 3893 12357 3927
rect 12391 3924 12403 3927
rect 12452 3924 12480 4091
rect 12544 4004 12572 4091
rect 12894 4088 12900 4140
rect 12952 4088 12958 4140
rect 13722 4088 13728 4140
rect 13780 4088 13786 4140
rect 13998 4088 14004 4140
rect 14056 4088 14062 4140
rect 14090 4088 14096 4140
rect 14148 4088 14154 4140
rect 14277 4131 14335 4137
rect 14277 4097 14289 4131
rect 14323 4097 14335 4131
rect 14277 4091 14335 4097
rect 14461 4131 14519 4137
rect 14461 4097 14473 4131
rect 14507 4128 14519 4131
rect 14734 4128 14740 4140
rect 14507 4100 14740 4128
rect 14507 4097 14519 4100
rect 14461 4091 14519 4097
rect 13541 4063 13599 4069
rect 13541 4029 13553 4063
rect 13587 4029 13599 4063
rect 13541 4023 13599 4029
rect 13909 4063 13967 4069
rect 13909 4029 13921 4063
rect 13955 4060 13967 4063
rect 14292 4060 14320 4091
rect 14734 4088 14740 4100
rect 14792 4088 14798 4140
rect 13955 4032 14320 4060
rect 13955 4029 13967 4032
rect 13909 4023 13967 4029
rect 12526 3952 12532 4004
rect 12584 3952 12590 4004
rect 13556 3936 13584 4023
rect 12618 3924 12624 3936
rect 12391 3896 12624 3924
rect 12391 3893 12403 3896
rect 12345 3887 12403 3893
rect 12618 3884 12624 3896
rect 12676 3884 12682 3936
rect 13538 3884 13544 3936
rect 13596 3884 13602 3936
rect 1104 3834 16376 3856
rect 1104 3782 2859 3834
rect 2911 3782 2923 3834
rect 2975 3782 2987 3834
rect 3039 3782 3051 3834
rect 3103 3782 3115 3834
rect 3167 3782 6677 3834
rect 6729 3782 6741 3834
rect 6793 3782 6805 3834
rect 6857 3782 6869 3834
rect 6921 3782 6933 3834
rect 6985 3782 10495 3834
rect 10547 3782 10559 3834
rect 10611 3782 10623 3834
rect 10675 3782 10687 3834
rect 10739 3782 10751 3834
rect 10803 3782 14313 3834
rect 14365 3782 14377 3834
rect 14429 3782 14441 3834
rect 14493 3782 14505 3834
rect 14557 3782 14569 3834
rect 14621 3782 16376 3834
rect 1104 3760 16376 3782
rect 5350 3680 5356 3732
rect 5408 3720 5414 3732
rect 6270 3720 6276 3732
rect 5408 3692 6276 3720
rect 5408 3680 5414 3692
rect 6270 3680 6276 3692
rect 6328 3680 6334 3732
rect 6365 3723 6423 3729
rect 6365 3689 6377 3723
rect 6411 3720 6423 3723
rect 7006 3720 7012 3732
rect 6411 3692 7012 3720
rect 6411 3689 6423 3692
rect 6365 3683 6423 3689
rect 7006 3680 7012 3692
rect 7064 3680 7070 3732
rect 7834 3680 7840 3732
rect 7892 3680 7898 3732
rect 8294 3680 8300 3732
rect 8352 3680 8358 3732
rect 9122 3680 9128 3732
rect 9180 3720 9186 3732
rect 9401 3723 9459 3729
rect 9401 3720 9413 3723
rect 9180 3692 9413 3720
rect 9180 3680 9186 3692
rect 9401 3689 9413 3692
rect 9447 3689 9459 3723
rect 9401 3683 9459 3689
rect 9674 3680 9680 3732
rect 9732 3680 9738 3732
rect 13722 3680 13728 3732
rect 13780 3680 13786 3732
rect 13909 3723 13967 3729
rect 13909 3689 13921 3723
rect 13955 3720 13967 3723
rect 13998 3720 14004 3732
rect 13955 3692 14004 3720
rect 13955 3689 13967 3692
rect 13909 3683 13967 3689
rect 13998 3680 14004 3692
rect 14056 3680 14062 3732
rect 5828 3624 6684 3652
rect 1673 3587 1731 3593
rect 1673 3553 1685 3587
rect 1719 3584 1731 3587
rect 3418 3584 3424 3596
rect 1719 3556 3424 3584
rect 1719 3553 1731 3556
rect 1673 3547 1731 3553
rect 3418 3544 3424 3556
rect 3476 3544 3482 3596
rect 4430 3544 4436 3596
rect 4488 3584 4494 3596
rect 5828 3584 5856 3624
rect 4488 3556 5856 3584
rect 4488 3544 4494 3556
rect 934 3476 940 3528
rect 992 3516 998 3528
rect 5828 3525 5856 3556
rect 6086 3544 6092 3596
rect 6144 3544 6150 3596
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 992 3488 1409 3516
rect 992 3476 998 3488
rect 1397 3485 1409 3488
rect 1443 3485 1455 3519
rect 1397 3479 1455 3485
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3485 4399 3519
rect 4341 3479 4399 3485
rect 5813 3519 5871 3525
rect 5813 3485 5825 3519
rect 5859 3485 5871 3519
rect 5813 3479 5871 3485
rect 5905 3519 5963 3525
rect 5905 3485 5917 3519
rect 5951 3485 5963 3519
rect 6104 3516 6132 3544
rect 6181 3519 6239 3525
rect 6181 3516 6193 3519
rect 6104 3488 6193 3516
rect 5905 3479 5963 3485
rect 6181 3485 6193 3488
rect 6227 3485 6239 3519
rect 6181 3479 6239 3485
rect 4356 3448 4384 3479
rect 4614 3448 4620 3460
rect 4356 3420 4620 3448
rect 4614 3408 4620 3420
rect 4672 3408 4678 3460
rect 5920 3448 5948 3479
rect 6270 3476 6276 3528
rect 6328 3516 6334 3528
rect 6656 3525 6684 3624
rect 6730 3612 6736 3664
rect 6788 3612 6794 3664
rect 6914 3612 6920 3664
rect 6972 3652 6978 3664
rect 7852 3652 7880 3680
rect 6972 3624 7880 3652
rect 8312 3652 8340 3680
rect 8312 3624 9536 3652
rect 6972 3612 6978 3624
rect 6457 3519 6515 3525
rect 6457 3516 6469 3519
rect 6328 3488 6469 3516
rect 6328 3476 6334 3488
rect 6457 3485 6469 3488
rect 6503 3485 6515 3519
rect 6457 3479 6515 3485
rect 6641 3519 6699 3525
rect 6641 3485 6653 3519
rect 6687 3516 6699 3519
rect 6733 3519 6791 3525
rect 6733 3516 6745 3519
rect 6687 3488 6745 3516
rect 6687 3485 6699 3488
rect 6641 3479 6699 3485
rect 6733 3485 6745 3488
rect 6779 3485 6791 3519
rect 6733 3479 6791 3485
rect 6917 3519 6975 3525
rect 6917 3485 6929 3519
rect 6963 3485 6975 3519
rect 6917 3479 6975 3485
rect 8113 3519 8171 3525
rect 8113 3485 8125 3519
rect 8159 3516 8171 3519
rect 8202 3516 8208 3528
rect 8159 3488 8208 3516
rect 8159 3485 8171 3488
rect 8113 3479 8171 3485
rect 6362 3448 6368 3460
rect 5920 3420 6368 3448
rect 6362 3408 6368 3420
rect 6420 3408 6426 3460
rect 4154 3340 4160 3392
rect 4212 3340 4218 3392
rect 5626 3340 5632 3392
rect 5684 3340 5690 3392
rect 5810 3340 5816 3392
rect 5868 3380 5874 3392
rect 5997 3383 6055 3389
rect 5997 3380 6009 3383
rect 5868 3352 6009 3380
rect 5868 3340 5874 3352
rect 5997 3349 6009 3352
rect 6043 3349 6055 3383
rect 6472 3380 6500 3479
rect 6546 3408 6552 3460
rect 6604 3408 6610 3460
rect 6932 3380 6960 3479
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3485 9367 3519
rect 9508 3516 9536 3624
rect 9585 3587 9643 3593
rect 9585 3553 9597 3587
rect 9631 3584 9643 3587
rect 9692 3584 9720 3680
rect 9631 3556 9720 3584
rect 9784 3624 13032 3652
rect 9631 3553 9643 3556
rect 9585 3547 9643 3553
rect 9784 3516 9812 3624
rect 12618 3544 12624 3596
rect 12676 3544 12682 3596
rect 12526 3516 12532 3528
rect 9508 3488 9812 3516
rect 12406 3488 12532 3516
rect 9309 3479 9367 3485
rect 9324 3392 9352 3479
rect 9585 3451 9643 3457
rect 9585 3417 9597 3451
rect 9631 3448 9643 3451
rect 12406 3448 12434 3488
rect 12526 3476 12532 3488
rect 12584 3516 12590 3528
rect 12713 3519 12771 3525
rect 12713 3516 12725 3519
rect 12584 3488 12725 3516
rect 12584 3476 12590 3488
rect 12713 3485 12725 3488
rect 12759 3485 12771 3519
rect 13004 3516 13032 3624
rect 13081 3587 13139 3593
rect 13081 3553 13093 3587
rect 13127 3584 13139 3587
rect 13633 3587 13691 3593
rect 13633 3584 13645 3587
rect 13127 3556 13645 3584
rect 13127 3553 13139 3556
rect 13081 3547 13139 3553
rect 13633 3553 13645 3556
rect 13679 3584 13691 3587
rect 13740 3584 13768 3680
rect 13679 3556 13768 3584
rect 14016 3584 14044 3680
rect 15930 3612 15936 3664
rect 15988 3612 15994 3664
rect 14185 3587 14243 3593
rect 14185 3584 14197 3587
rect 14016 3556 14197 3584
rect 13679 3553 13691 3556
rect 13633 3547 13691 3553
rect 14185 3553 14197 3556
rect 14231 3553 14243 3587
rect 14185 3547 14243 3553
rect 14645 3587 14703 3593
rect 14645 3553 14657 3587
rect 14691 3553 14703 3587
rect 14645 3547 14703 3553
rect 13538 3516 13544 3528
rect 13004 3488 13544 3516
rect 12713 3479 12771 3485
rect 13538 3476 13544 3488
rect 13596 3476 13602 3528
rect 14277 3519 14335 3525
rect 14277 3485 14289 3519
rect 14323 3485 14335 3519
rect 14660 3516 14688 3547
rect 15749 3519 15807 3525
rect 15749 3516 15761 3519
rect 14660 3488 15761 3516
rect 14277 3479 14335 3485
rect 15749 3485 15761 3488
rect 15795 3485 15807 3519
rect 15749 3479 15807 3485
rect 14090 3448 14096 3460
rect 9631 3420 12434 3448
rect 13188 3420 14096 3448
rect 9631 3417 9643 3420
rect 9585 3411 9643 3417
rect 13188 3392 13216 3420
rect 14090 3408 14096 3420
rect 14148 3448 14154 3460
rect 14292 3448 14320 3479
rect 14148 3420 14320 3448
rect 14148 3408 14154 3420
rect 6472 3352 6960 3380
rect 5997 3343 6055 3349
rect 7006 3340 7012 3392
rect 7064 3380 7070 3392
rect 7929 3383 7987 3389
rect 7929 3380 7941 3383
rect 7064 3352 7941 3380
rect 7064 3340 7070 3352
rect 7929 3349 7941 3352
rect 7975 3349 7987 3383
rect 7929 3343 7987 3349
rect 9306 3340 9312 3392
rect 9364 3340 9370 3392
rect 13170 3340 13176 3392
rect 13228 3340 13234 3392
rect 1104 3290 16376 3312
rect 1104 3238 3519 3290
rect 3571 3238 3583 3290
rect 3635 3238 3647 3290
rect 3699 3238 3711 3290
rect 3763 3238 3775 3290
rect 3827 3238 7337 3290
rect 7389 3238 7401 3290
rect 7453 3238 7465 3290
rect 7517 3238 7529 3290
rect 7581 3238 7593 3290
rect 7645 3238 11155 3290
rect 11207 3238 11219 3290
rect 11271 3238 11283 3290
rect 11335 3238 11347 3290
rect 11399 3238 11411 3290
rect 11463 3238 14973 3290
rect 15025 3238 15037 3290
rect 15089 3238 15101 3290
rect 15153 3238 15165 3290
rect 15217 3238 15229 3290
rect 15281 3238 16376 3290
rect 1104 3216 16376 3238
rect 3326 3136 3332 3188
rect 3384 3136 3390 3188
rect 4154 3136 4160 3188
rect 4212 3136 4218 3188
rect 4249 3179 4307 3185
rect 4249 3145 4261 3179
rect 4295 3176 4307 3179
rect 4614 3176 4620 3188
rect 4295 3148 4620 3176
rect 4295 3145 4307 3148
rect 4249 3139 4307 3145
rect 4614 3136 4620 3148
rect 4672 3136 4678 3188
rect 5626 3136 5632 3188
rect 5684 3136 5690 3188
rect 6181 3179 6239 3185
rect 6181 3145 6193 3179
rect 6227 3145 6239 3179
rect 6181 3139 6239 3145
rect 934 3000 940 3052
rect 992 3040 998 3052
rect 1397 3043 1455 3049
rect 1397 3040 1409 3043
rect 992 3012 1409 3040
rect 992 3000 998 3012
rect 1397 3009 1409 3012
rect 1443 3009 1455 3043
rect 1397 3003 1455 3009
rect 2961 3043 3019 3049
rect 2961 3009 2973 3043
rect 3007 3040 3019 3043
rect 3344 3040 3372 3136
rect 4172 3108 4200 3136
rect 3712 3080 4200 3108
rect 3712 3049 3740 3080
rect 3007 3012 3372 3040
rect 3007 3009 3019 3012
rect 2961 3003 3019 3009
rect 1946 2932 1952 2984
rect 2004 2932 2010 2984
rect 3344 2904 3372 3012
rect 3697 3043 3755 3049
rect 3697 3009 3709 3043
rect 3743 3009 3755 3043
rect 4157 3043 4215 3049
rect 4157 3040 4169 3043
rect 3697 3003 3755 3009
rect 3804 3012 4169 3040
rect 3421 2975 3479 2981
rect 3421 2941 3433 2975
rect 3467 2972 3479 2975
rect 3605 2975 3663 2981
rect 3605 2972 3617 2975
rect 3467 2944 3617 2972
rect 3467 2941 3479 2944
rect 3421 2935 3479 2941
rect 3605 2941 3617 2944
rect 3651 2941 3663 2975
rect 3605 2935 3663 2941
rect 3804 2904 3832 3012
rect 4157 3009 4169 3012
rect 4203 3009 4215 3043
rect 4157 3003 4215 3009
rect 4433 3043 4491 3049
rect 4433 3009 4445 3043
rect 4479 3009 4491 3043
rect 4433 3003 4491 3009
rect 5169 3043 5227 3049
rect 5169 3009 5181 3043
rect 5215 3040 5227 3043
rect 5350 3040 5356 3052
rect 5215 3012 5356 3040
rect 5215 3009 5227 3012
rect 5169 3003 5227 3009
rect 3970 2932 3976 2984
rect 4028 2972 4034 2984
rect 4448 2972 4476 3003
rect 5350 3000 5356 3012
rect 5408 3000 5414 3052
rect 4028 2944 4476 2972
rect 5261 2975 5319 2981
rect 4028 2932 4034 2944
rect 5261 2941 5273 2975
rect 5307 2972 5319 2975
rect 5644 2972 5672 3136
rect 6196 3108 6224 3139
rect 7006 3136 7012 3188
rect 7064 3136 7070 3188
rect 8313 3179 8371 3185
rect 8313 3176 8325 3179
rect 7208 3148 8325 3176
rect 7208 3117 7236 3148
rect 8313 3145 8325 3148
rect 8359 3145 8371 3179
rect 8570 3176 8576 3188
rect 8313 3139 8371 3145
rect 8404 3148 8576 3176
rect 7193 3111 7251 3117
rect 7193 3108 7205 3111
rect 6196 3080 7205 3108
rect 7193 3077 7205 3080
rect 7239 3077 7251 3111
rect 7193 3071 7251 3077
rect 7377 3111 7435 3117
rect 7377 3077 7389 3111
rect 7423 3108 7435 3111
rect 7650 3108 7656 3120
rect 7423 3080 7656 3108
rect 7423 3077 7435 3080
rect 7377 3071 7435 3077
rect 7650 3068 7656 3080
rect 7708 3068 7714 3120
rect 7853 3111 7911 3117
rect 7853 3108 7865 3111
rect 7760 3080 7865 3108
rect 5810 3000 5816 3052
rect 5868 3000 5874 3052
rect 6914 3000 6920 3052
rect 6972 3000 6978 3052
rect 7285 3043 7343 3049
rect 7285 3009 7297 3043
rect 7331 3040 7343 3043
rect 7561 3043 7619 3049
rect 7331 3012 7420 3040
rect 7331 3009 7343 3012
rect 7285 3003 7343 3009
rect 5307 2944 5672 2972
rect 5721 2975 5779 2981
rect 5307 2941 5319 2944
rect 5261 2935 5319 2941
rect 5721 2941 5733 2975
rect 5767 2941 5779 2975
rect 5721 2935 5779 2941
rect 3344 2876 3832 2904
rect 3237 2839 3295 2845
rect 3237 2805 3249 2839
rect 3283 2836 3295 2839
rect 3988 2836 4016 2932
rect 4065 2907 4123 2913
rect 4065 2873 4077 2907
rect 4111 2904 4123 2907
rect 4338 2904 4344 2916
rect 4111 2876 4344 2904
rect 4111 2873 4123 2876
rect 4065 2867 4123 2873
rect 4338 2864 4344 2876
rect 4396 2864 4402 2916
rect 5537 2907 5595 2913
rect 5537 2873 5549 2907
rect 5583 2904 5595 2907
rect 5736 2904 5764 2935
rect 5583 2876 5764 2904
rect 5583 2873 5595 2876
rect 5537 2867 5595 2873
rect 3283 2808 4016 2836
rect 4617 2839 4675 2845
rect 3283 2805 3295 2808
rect 3237 2799 3295 2805
rect 4617 2805 4629 2839
rect 4663 2836 4675 2839
rect 5828 2836 5856 3000
rect 7190 2932 7196 2984
rect 7248 2972 7254 2984
rect 7392 2972 7420 3012
rect 7561 3009 7573 3043
rect 7607 3040 7619 3043
rect 7760 3040 7788 3080
rect 7853 3077 7865 3080
rect 7899 3077 7911 3111
rect 7853 3071 7911 3077
rect 8113 3111 8171 3117
rect 8113 3077 8125 3111
rect 8159 3108 8171 3111
rect 8202 3108 8208 3120
rect 8159 3080 8208 3108
rect 8159 3077 8171 3080
rect 8113 3071 8171 3077
rect 8202 3068 8208 3080
rect 8260 3068 8266 3120
rect 8404 3108 8432 3148
rect 8570 3136 8576 3148
rect 8628 3136 8634 3188
rect 12069 3179 12127 3185
rect 8772 3148 11652 3176
rect 8328 3080 8432 3108
rect 8328 3040 8356 3080
rect 8478 3068 8484 3120
rect 8536 3108 8542 3120
rect 8772 3108 8800 3148
rect 8536 3080 8800 3108
rect 8536 3068 8542 3080
rect 7607 3012 7788 3040
rect 7607 3009 7619 3012
rect 7561 3003 7619 3009
rect 7760 2984 7788 3012
rect 7944 3012 8356 3040
rect 7248 2944 7420 2972
rect 7248 2932 7254 2944
rect 4663 2808 5856 2836
rect 4663 2805 4675 2808
rect 4617 2799 4675 2805
rect 7190 2796 7196 2848
rect 7248 2796 7254 2848
rect 7392 2836 7420 2944
rect 7742 2932 7748 2984
rect 7800 2932 7806 2984
rect 7561 2907 7619 2913
rect 7561 2873 7573 2907
rect 7607 2904 7619 2907
rect 7944 2904 7972 3012
rect 8570 3000 8576 3052
rect 8628 3000 8634 3052
rect 8772 3049 8800 3080
rect 9306 3068 9312 3120
rect 9364 3068 9370 3120
rect 8757 3043 8815 3049
rect 8757 3009 8769 3043
rect 8803 3009 8815 3043
rect 8757 3003 8815 3009
rect 8849 3043 8907 3049
rect 8849 3009 8861 3043
rect 8895 3009 8907 3043
rect 8849 3003 8907 3009
rect 8941 3043 8999 3049
rect 8941 3009 8953 3043
rect 8987 3040 8999 3043
rect 9324 3040 9352 3068
rect 9401 3043 9459 3049
rect 9401 3040 9413 3043
rect 8987 3012 9413 3040
rect 8987 3009 8999 3012
rect 8941 3003 8999 3009
rect 9401 3009 9413 3012
rect 9447 3009 9459 3043
rect 9401 3003 9459 3009
rect 7607 2876 7972 2904
rect 8021 2907 8079 2913
rect 7607 2873 7619 2876
rect 7561 2867 7619 2873
rect 8021 2873 8033 2907
rect 8067 2904 8079 2907
rect 8386 2904 8392 2916
rect 8067 2876 8392 2904
rect 8067 2873 8079 2876
rect 8021 2867 8079 2873
rect 8386 2864 8392 2876
rect 8444 2864 8450 2916
rect 8864 2904 8892 3003
rect 9766 3000 9772 3052
rect 9824 3040 9830 3052
rect 10229 3043 10287 3049
rect 10229 3040 10241 3043
rect 9824 3012 10241 3040
rect 9824 3000 9830 3012
rect 10229 3009 10241 3012
rect 10275 3009 10287 3043
rect 10229 3003 10287 3009
rect 11149 3043 11207 3049
rect 11149 3009 11161 3043
rect 11195 3009 11207 3043
rect 11149 3003 11207 3009
rect 11333 3043 11391 3049
rect 11333 3009 11345 3043
rect 11379 3040 11391 3043
rect 11624 3040 11652 3148
rect 12069 3145 12081 3179
rect 12115 3176 12127 3179
rect 12115 3148 12434 3176
rect 12115 3145 12127 3148
rect 12069 3139 12127 3145
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 11379 3012 11560 3040
rect 11624 3012 11713 3040
rect 11379 3009 11391 3012
rect 11333 3003 11391 3009
rect 9122 2932 9128 2984
rect 9180 2972 9186 2984
rect 9309 2975 9367 2981
rect 9309 2972 9321 2975
rect 9180 2944 9321 2972
rect 9180 2932 9186 2944
rect 9309 2941 9321 2944
rect 9355 2941 9367 2975
rect 9309 2935 9367 2941
rect 10321 2975 10379 2981
rect 10321 2941 10333 2975
rect 10367 2972 10379 2975
rect 10410 2972 10416 2984
rect 10367 2944 10416 2972
rect 10367 2941 10379 2944
rect 10321 2935 10379 2941
rect 8496 2876 8892 2904
rect 9769 2907 9827 2913
rect 8496 2848 8524 2876
rect 9769 2873 9781 2907
rect 9815 2904 9827 2907
rect 10336 2904 10364 2935
rect 10410 2932 10416 2944
rect 10468 2932 10474 2984
rect 9815 2876 10364 2904
rect 10597 2907 10655 2913
rect 9815 2873 9827 2876
rect 9769 2867 9827 2873
rect 10597 2873 10609 2907
rect 10643 2904 10655 2907
rect 11164 2904 11192 3003
rect 11422 2932 11428 2984
rect 11480 2932 11486 2984
rect 11440 2904 11468 2932
rect 10643 2876 11468 2904
rect 11532 2904 11560 3012
rect 11701 3009 11713 3012
rect 11747 3040 11759 3043
rect 12161 3043 12219 3049
rect 12161 3040 12173 3043
rect 11747 3012 12173 3040
rect 11747 3009 11759 3012
rect 11701 3003 11759 3009
rect 12161 3009 12173 3012
rect 12207 3009 12219 3043
rect 12161 3003 12219 3009
rect 11606 2932 11612 2984
rect 11664 2932 11670 2984
rect 12406 2916 12434 3148
rect 12253 2907 12311 2913
rect 12253 2904 12265 2907
rect 11532 2876 12265 2904
rect 10643 2873 10655 2876
rect 10597 2867 10655 2873
rect 12253 2873 12265 2876
rect 12299 2873 12311 2907
rect 12406 2876 12440 2916
rect 12253 2867 12311 2873
rect 12434 2864 12440 2876
rect 12492 2864 12498 2916
rect 7837 2839 7895 2845
rect 7837 2836 7849 2839
rect 7392 2808 7849 2836
rect 7837 2805 7849 2808
rect 7883 2805 7895 2839
rect 7837 2799 7895 2805
rect 7926 2796 7932 2848
rect 7984 2836 7990 2848
rect 8297 2839 8355 2845
rect 8297 2836 8309 2839
rect 7984 2808 8309 2836
rect 7984 2796 7990 2808
rect 8297 2805 8309 2808
rect 8343 2805 8355 2839
rect 8297 2799 8355 2805
rect 8478 2796 8484 2848
rect 8536 2796 8542 2848
rect 8570 2796 8576 2848
rect 8628 2796 8634 2848
rect 10870 2796 10876 2848
rect 10928 2796 10934 2848
rect 11149 2839 11207 2845
rect 11149 2805 11161 2839
rect 11195 2836 11207 2839
rect 13170 2836 13176 2848
rect 11195 2808 13176 2836
rect 11195 2805 11207 2808
rect 11149 2799 11207 2805
rect 13170 2796 13176 2808
rect 13228 2796 13234 2848
rect 1104 2746 16376 2768
rect 1104 2694 2859 2746
rect 2911 2694 2923 2746
rect 2975 2694 2987 2746
rect 3039 2694 3051 2746
rect 3103 2694 3115 2746
rect 3167 2694 6677 2746
rect 6729 2694 6741 2746
rect 6793 2694 6805 2746
rect 6857 2694 6869 2746
rect 6921 2694 6933 2746
rect 6985 2694 10495 2746
rect 10547 2694 10559 2746
rect 10611 2694 10623 2746
rect 10675 2694 10687 2746
rect 10739 2694 10751 2746
rect 10803 2694 14313 2746
rect 14365 2694 14377 2746
rect 14429 2694 14441 2746
rect 14493 2694 14505 2746
rect 14557 2694 14569 2746
rect 14621 2694 16376 2746
rect 1104 2672 16376 2694
rect 7098 2592 7104 2644
rect 7156 2632 7162 2644
rect 7377 2635 7435 2641
rect 7377 2632 7389 2635
rect 7156 2604 7389 2632
rect 7156 2592 7162 2604
rect 7377 2601 7389 2604
rect 7423 2601 7435 2635
rect 7377 2595 7435 2601
rect 7742 2592 7748 2644
rect 7800 2592 7806 2644
rect 8018 2592 8024 2644
rect 8076 2592 8082 2644
rect 9309 2635 9367 2641
rect 9309 2601 9321 2635
rect 9355 2632 9367 2635
rect 9398 2632 9404 2644
rect 9355 2604 9404 2632
rect 9355 2601 9367 2604
rect 9309 2595 9367 2601
rect 9398 2592 9404 2604
rect 9456 2592 9462 2644
rect 10505 2635 10563 2641
rect 10505 2601 10517 2635
rect 10551 2632 10563 2635
rect 10870 2632 10876 2644
rect 10551 2604 10876 2632
rect 10551 2601 10563 2604
rect 10505 2595 10563 2601
rect 10870 2592 10876 2604
rect 10928 2592 10934 2644
rect 7190 2524 7196 2576
rect 7248 2524 7254 2576
rect 7208 2496 7236 2524
rect 8478 2496 8484 2508
rect 7208 2468 7788 2496
rect 4338 2388 4344 2440
rect 4396 2428 4402 2440
rect 4709 2431 4767 2437
rect 4709 2428 4721 2431
rect 4396 2400 4721 2428
rect 4396 2388 4402 2400
rect 4709 2397 4721 2400
rect 4755 2397 4767 2431
rect 4709 2391 4767 2397
rect 7190 2388 7196 2440
rect 7248 2388 7254 2440
rect 7760 2437 7788 2468
rect 7944 2468 8484 2496
rect 7944 2437 7972 2468
rect 8478 2456 8484 2468
rect 8536 2456 8542 2508
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2397 7803 2431
rect 7745 2391 7803 2397
rect 7929 2431 7987 2437
rect 7929 2397 7941 2431
rect 7975 2397 7987 2431
rect 7929 2391 7987 2397
rect 8205 2431 8263 2437
rect 8205 2397 8217 2431
rect 8251 2397 8263 2431
rect 8205 2391 8263 2397
rect 8220 2360 8248 2391
rect 8570 2388 8576 2440
rect 8628 2428 8634 2440
rect 8665 2431 8723 2437
rect 8665 2428 8677 2431
rect 8628 2400 8677 2428
rect 8628 2388 8634 2400
rect 8665 2397 8677 2400
rect 8711 2397 8723 2431
rect 8665 2391 8723 2397
rect 9122 2388 9128 2440
rect 9180 2388 9186 2440
rect 9950 2388 9956 2440
rect 10008 2428 10014 2440
rect 10321 2431 10379 2437
rect 10321 2428 10333 2431
rect 10008 2400 10333 2428
rect 10008 2388 10014 2400
rect 10321 2397 10333 2400
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 10410 2388 10416 2440
rect 10468 2428 10474 2440
rect 10505 2431 10563 2437
rect 10505 2428 10517 2431
rect 10468 2400 10517 2428
rect 10468 2388 10474 2400
rect 10505 2397 10517 2400
rect 10551 2397 10563 2431
rect 10505 2391 10563 2397
rect 12434 2388 12440 2440
rect 12492 2388 12498 2440
rect 7760 2332 8248 2360
rect 7760 2304 7788 2332
rect 4522 2252 4528 2304
rect 4580 2292 4586 2304
rect 4801 2295 4859 2301
rect 4801 2292 4813 2295
rect 4580 2264 4813 2292
rect 4580 2252 4586 2264
rect 4801 2261 4813 2264
rect 4847 2261 4859 2295
rect 4801 2255 4859 2261
rect 7742 2252 7748 2304
rect 7800 2252 7806 2304
rect 8386 2252 8392 2304
rect 8444 2252 8450 2304
rect 12342 2252 12348 2304
rect 12400 2292 12406 2304
rect 12529 2295 12587 2301
rect 12529 2292 12541 2295
rect 12400 2264 12541 2292
rect 12400 2252 12406 2264
rect 12529 2261 12541 2264
rect 12575 2261 12587 2295
rect 12529 2255 12587 2261
rect 1104 2202 16376 2224
rect 1104 2150 3519 2202
rect 3571 2150 3583 2202
rect 3635 2150 3647 2202
rect 3699 2150 3711 2202
rect 3763 2150 3775 2202
rect 3827 2150 7337 2202
rect 7389 2150 7401 2202
rect 7453 2150 7465 2202
rect 7517 2150 7529 2202
rect 7581 2150 7593 2202
rect 7645 2150 11155 2202
rect 11207 2150 11219 2202
rect 11271 2150 11283 2202
rect 11335 2150 11347 2202
rect 11399 2150 11411 2202
rect 11463 2150 14973 2202
rect 15025 2150 15037 2202
rect 15089 2150 15101 2202
rect 15153 2150 15165 2202
rect 15217 2150 15229 2202
rect 15281 2150 16376 2202
rect 1104 2128 16376 2150
<< via1 >>
rect 3519 17382 3571 17434
rect 3583 17382 3635 17434
rect 3647 17382 3699 17434
rect 3711 17382 3763 17434
rect 3775 17382 3827 17434
rect 7337 17382 7389 17434
rect 7401 17382 7453 17434
rect 7465 17382 7517 17434
rect 7529 17382 7581 17434
rect 7593 17382 7645 17434
rect 11155 17382 11207 17434
rect 11219 17382 11271 17434
rect 11283 17382 11335 17434
rect 11347 17382 11399 17434
rect 11411 17382 11463 17434
rect 14973 17382 15025 17434
rect 15037 17382 15089 17434
rect 15101 17382 15153 17434
rect 15165 17382 15217 17434
rect 15229 17382 15281 17434
rect 13820 17280 13872 17332
rect 14832 17280 14884 17332
rect 12440 17212 12492 17264
rect 7196 17187 7248 17196
rect 7196 17153 7205 17187
rect 7205 17153 7239 17187
rect 7239 17153 7248 17187
rect 7196 17144 7248 17153
rect 7288 17144 7340 17196
rect 8024 17144 8076 17196
rect 10324 17187 10376 17196
rect 10324 17153 10333 17187
rect 10333 17153 10367 17187
rect 10367 17153 10376 17187
rect 10324 17144 10376 17153
rect 10416 17187 10468 17196
rect 10416 17153 10425 17187
rect 10425 17153 10459 17187
rect 10459 17153 10468 17187
rect 10416 17144 10468 17153
rect 9864 17076 9916 17128
rect 12164 17187 12216 17196
rect 12164 17153 12173 17187
rect 12173 17153 12207 17187
rect 12207 17153 12216 17187
rect 12164 17144 12216 17153
rect 12808 17144 12860 17196
rect 10876 17076 10928 17128
rect 12072 17076 12124 17128
rect 14188 17187 14240 17196
rect 14188 17153 14197 17187
rect 14197 17153 14231 17187
rect 14231 17153 14240 17187
rect 14188 17144 14240 17153
rect 15016 17187 15068 17196
rect 15016 17153 15025 17187
rect 15025 17153 15059 17187
rect 15059 17153 15068 17187
rect 15016 17144 15068 17153
rect 7472 17008 7524 17060
rect 12624 17008 12676 17060
rect 9036 16940 9088 16992
rect 11612 16940 11664 16992
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 12900 16940 12952 16949
rect 2859 16838 2911 16890
rect 2923 16838 2975 16890
rect 2987 16838 3039 16890
rect 3051 16838 3103 16890
rect 3115 16838 3167 16890
rect 6677 16838 6729 16890
rect 6741 16838 6793 16890
rect 6805 16838 6857 16890
rect 6869 16838 6921 16890
rect 6933 16838 6985 16890
rect 10495 16838 10547 16890
rect 10559 16838 10611 16890
rect 10623 16838 10675 16890
rect 10687 16838 10739 16890
rect 10751 16838 10803 16890
rect 14313 16838 14365 16890
rect 14377 16838 14429 16890
rect 14441 16838 14493 16890
rect 14505 16838 14557 16890
rect 14569 16838 14621 16890
rect 7196 16736 7248 16788
rect 7472 16736 7524 16788
rect 8024 16736 8076 16788
rect 6000 16532 6052 16584
rect 7196 16532 7248 16584
rect 8208 16600 8260 16652
rect 6552 16464 6604 16516
rect 7932 16575 7984 16584
rect 7932 16541 7941 16575
rect 7941 16541 7975 16575
rect 7975 16541 7984 16575
rect 7932 16532 7984 16541
rect 8024 16575 8076 16584
rect 8024 16541 8033 16575
rect 8033 16541 8067 16575
rect 8067 16541 8076 16575
rect 8024 16532 8076 16541
rect 9036 16736 9088 16788
rect 10140 16736 10192 16788
rect 10416 16736 10468 16788
rect 10508 16736 10560 16788
rect 8944 16532 8996 16584
rect 10232 16575 10284 16584
rect 10232 16541 10241 16575
rect 10241 16541 10275 16575
rect 10275 16541 10284 16575
rect 10232 16532 10284 16541
rect 10324 16575 10376 16584
rect 10324 16541 10333 16575
rect 10333 16541 10367 16575
rect 10367 16541 10376 16575
rect 10324 16532 10376 16541
rect 12072 16779 12124 16788
rect 12072 16745 12081 16779
rect 12081 16745 12115 16779
rect 12115 16745 12124 16779
rect 12072 16736 12124 16745
rect 12164 16779 12216 16788
rect 12164 16745 12173 16779
rect 12173 16745 12207 16779
rect 12207 16745 12216 16779
rect 12164 16736 12216 16745
rect 14188 16736 14240 16788
rect 15016 16736 15068 16788
rect 12532 16668 12584 16720
rect 12900 16643 12952 16652
rect 6460 16439 6512 16448
rect 6460 16405 6469 16439
rect 6469 16405 6503 16439
rect 6503 16405 6512 16439
rect 6460 16396 6512 16405
rect 7748 16396 7800 16448
rect 9864 16396 9916 16448
rect 12900 16609 12909 16643
rect 12909 16609 12943 16643
rect 12943 16609 12952 16643
rect 12900 16600 12952 16609
rect 14372 16643 14424 16652
rect 14372 16609 14381 16643
rect 14381 16609 14415 16643
rect 14415 16609 14424 16643
rect 14372 16600 14424 16609
rect 10876 16507 10928 16516
rect 10876 16473 10901 16507
rect 10901 16473 10928 16507
rect 10876 16464 10928 16473
rect 12624 16575 12676 16584
rect 12624 16541 12633 16575
rect 12633 16541 12667 16575
rect 12667 16541 12676 16575
rect 12624 16532 12676 16541
rect 12716 16575 12768 16584
rect 12716 16541 12725 16575
rect 12725 16541 12759 16575
rect 12759 16541 12768 16575
rect 12716 16532 12768 16541
rect 11060 16439 11112 16448
rect 11060 16405 11069 16439
rect 11069 16405 11103 16439
rect 11103 16405 11112 16439
rect 11060 16396 11112 16405
rect 11888 16439 11940 16448
rect 11888 16405 11913 16439
rect 11913 16405 11940 16439
rect 13728 16532 13780 16584
rect 11888 16396 11940 16405
rect 12900 16396 12952 16448
rect 13636 16396 13688 16448
rect 3519 16294 3571 16346
rect 3583 16294 3635 16346
rect 3647 16294 3699 16346
rect 3711 16294 3763 16346
rect 3775 16294 3827 16346
rect 7337 16294 7389 16346
rect 7401 16294 7453 16346
rect 7465 16294 7517 16346
rect 7529 16294 7581 16346
rect 7593 16294 7645 16346
rect 11155 16294 11207 16346
rect 11219 16294 11271 16346
rect 11283 16294 11335 16346
rect 11347 16294 11399 16346
rect 11411 16294 11463 16346
rect 14973 16294 15025 16346
rect 15037 16294 15089 16346
rect 15101 16294 15153 16346
rect 15165 16294 15217 16346
rect 15229 16294 15281 16346
rect 7748 16192 7800 16244
rect 11888 16192 11940 16244
rect 4160 16056 4212 16108
rect 5632 16099 5684 16108
rect 5632 16065 5641 16099
rect 5641 16065 5675 16099
rect 5675 16065 5684 16099
rect 5632 16056 5684 16065
rect 6828 16056 6880 16108
rect 7104 16056 7156 16108
rect 7472 16167 7524 16176
rect 7472 16133 7497 16167
rect 7497 16133 7524 16167
rect 7472 16124 7524 16133
rect 8208 16124 8260 16176
rect 10324 16124 10376 16176
rect 12072 16124 12124 16176
rect 12716 16192 12768 16244
rect 12900 16192 12952 16244
rect 13636 16235 13688 16244
rect 13636 16201 13645 16235
rect 13645 16201 13679 16235
rect 13679 16201 13688 16235
rect 13636 16192 13688 16201
rect 11060 16056 11112 16108
rect 11612 16056 11664 16108
rect 12532 16056 12584 16108
rect 13728 16124 13780 16176
rect 13912 16124 13964 16176
rect 6000 15920 6052 15972
rect 6460 15920 6512 15972
rect 10232 15988 10284 16040
rect 10140 15963 10192 15972
rect 10140 15929 10149 15963
rect 10149 15929 10183 15963
rect 10183 15929 10192 15963
rect 10140 15920 10192 15929
rect 12808 15920 12860 15972
rect 14372 15963 14424 15972
rect 14372 15929 14381 15963
rect 14381 15929 14415 15963
rect 14415 15929 14424 15963
rect 14372 15920 14424 15929
rect 7748 15852 7800 15904
rect 7932 15852 7984 15904
rect 10416 15852 10468 15904
rect 13820 15895 13872 15904
rect 13820 15861 13829 15895
rect 13829 15861 13863 15895
rect 13863 15861 13872 15895
rect 13820 15852 13872 15861
rect 14188 15852 14240 15904
rect 2859 15750 2911 15802
rect 2923 15750 2975 15802
rect 2987 15750 3039 15802
rect 3051 15750 3103 15802
rect 3115 15750 3167 15802
rect 6677 15750 6729 15802
rect 6741 15750 6793 15802
rect 6805 15750 6857 15802
rect 6869 15750 6921 15802
rect 6933 15750 6985 15802
rect 10495 15750 10547 15802
rect 10559 15750 10611 15802
rect 10623 15750 10675 15802
rect 10687 15750 10739 15802
rect 10751 15750 10803 15802
rect 14313 15750 14365 15802
rect 14377 15750 14429 15802
rect 14441 15750 14493 15802
rect 14505 15750 14557 15802
rect 14569 15750 14621 15802
rect 6000 15648 6052 15700
rect 7196 15648 7248 15700
rect 7472 15648 7524 15700
rect 6460 15580 6512 15632
rect 9404 15580 9456 15632
rect 7012 15444 7064 15496
rect 7104 15444 7156 15496
rect 7196 15376 7248 15428
rect 6644 15308 6696 15360
rect 7012 15308 7064 15360
rect 9404 15308 9456 15360
rect 10324 15444 10376 15496
rect 14096 15376 14148 15428
rect 10232 15351 10284 15360
rect 10232 15317 10241 15351
rect 10241 15317 10275 15351
rect 10275 15317 10284 15351
rect 10232 15308 10284 15317
rect 12716 15308 12768 15360
rect 14188 15308 14240 15360
rect 16028 15308 16080 15360
rect 3519 15206 3571 15258
rect 3583 15206 3635 15258
rect 3647 15206 3699 15258
rect 3711 15206 3763 15258
rect 3775 15206 3827 15258
rect 7337 15206 7389 15258
rect 7401 15206 7453 15258
rect 7465 15206 7517 15258
rect 7529 15206 7581 15258
rect 7593 15206 7645 15258
rect 11155 15206 11207 15258
rect 11219 15206 11271 15258
rect 11283 15206 11335 15258
rect 11347 15206 11399 15258
rect 11411 15206 11463 15258
rect 14973 15206 15025 15258
rect 15037 15206 15089 15258
rect 15101 15206 15153 15258
rect 15165 15206 15217 15258
rect 15229 15206 15281 15258
rect 2136 14764 2188 14816
rect 3884 15036 3936 15088
rect 6552 15104 6604 15156
rect 2688 15011 2740 15020
rect 2688 14977 2697 15011
rect 2697 14977 2731 15011
rect 2731 14977 2740 15011
rect 2688 14968 2740 14977
rect 4160 14968 4212 15020
rect 4252 15011 4304 15020
rect 4252 14977 4261 15011
rect 4261 14977 4295 15011
rect 4295 14977 4304 15011
rect 4252 14968 4304 14977
rect 3792 14900 3844 14952
rect 5264 14968 5316 15020
rect 5632 14968 5684 15020
rect 7196 15036 7248 15088
rect 10232 15036 10284 15088
rect 7104 15011 7156 15020
rect 7104 14977 7113 15011
rect 7113 14977 7147 15011
rect 7147 14977 7156 15011
rect 7104 14968 7156 14977
rect 6552 14900 6604 14952
rect 7840 14900 7892 14952
rect 10600 14968 10652 15020
rect 12716 15036 12768 15088
rect 5172 14764 5224 14816
rect 7012 14764 7064 14816
rect 7196 14764 7248 14816
rect 10048 14764 10100 14816
rect 10140 14807 10192 14816
rect 10140 14773 10149 14807
rect 10149 14773 10183 14807
rect 10183 14773 10192 14807
rect 13912 14968 13964 15020
rect 13820 14943 13872 14952
rect 13820 14909 13829 14943
rect 13829 14909 13863 14943
rect 13863 14909 13872 14943
rect 14188 15011 14240 15020
rect 14188 14977 14197 15011
rect 14197 14977 14231 15011
rect 14231 14977 14240 15011
rect 14188 14968 14240 14977
rect 13820 14900 13872 14909
rect 14096 14943 14148 14952
rect 14096 14909 14105 14943
rect 14105 14909 14139 14943
rect 14139 14909 14148 14943
rect 14096 14900 14148 14909
rect 10140 14764 10192 14773
rect 10600 14764 10652 14816
rect 10968 14764 11020 14816
rect 12808 14764 12860 14816
rect 12992 14764 13044 14816
rect 2859 14662 2911 14714
rect 2923 14662 2975 14714
rect 2987 14662 3039 14714
rect 3051 14662 3103 14714
rect 3115 14662 3167 14714
rect 6677 14662 6729 14714
rect 6741 14662 6793 14714
rect 6805 14662 6857 14714
rect 6869 14662 6921 14714
rect 6933 14662 6985 14714
rect 10495 14662 10547 14714
rect 10559 14662 10611 14714
rect 10623 14662 10675 14714
rect 10687 14662 10739 14714
rect 10751 14662 10803 14714
rect 14313 14662 14365 14714
rect 14377 14662 14429 14714
rect 14441 14662 14493 14714
rect 14505 14662 14557 14714
rect 14569 14662 14621 14714
rect 4068 14560 4120 14612
rect 3332 14535 3384 14544
rect 3332 14501 3341 14535
rect 3341 14501 3375 14535
rect 3375 14501 3384 14535
rect 3332 14492 3384 14501
rect 940 14288 992 14340
rect 2596 14288 2648 14340
rect 2780 14331 2832 14340
rect 2780 14297 2789 14331
rect 2789 14297 2823 14331
rect 2823 14297 2832 14331
rect 2780 14288 2832 14297
rect 1400 14220 1452 14272
rect 2228 14220 2280 14272
rect 2688 14220 2740 14272
rect 3240 14356 3292 14408
rect 3516 14424 3568 14476
rect 3792 14467 3844 14476
rect 3792 14433 3801 14467
rect 3801 14433 3835 14467
rect 3835 14433 3844 14467
rect 3792 14424 3844 14433
rect 3884 14424 3936 14476
rect 4252 14467 4304 14476
rect 4252 14433 4262 14467
rect 4262 14433 4296 14467
rect 4296 14433 4304 14467
rect 5264 14560 5316 14612
rect 9404 14603 9456 14612
rect 9404 14569 9413 14603
rect 9413 14569 9447 14603
rect 9447 14569 9456 14603
rect 9404 14560 9456 14569
rect 10048 14603 10100 14612
rect 10048 14569 10057 14603
rect 10057 14569 10091 14603
rect 10091 14569 10100 14603
rect 10048 14560 10100 14569
rect 10968 14603 11020 14612
rect 10968 14569 10977 14603
rect 10977 14569 11011 14603
rect 11011 14569 11020 14603
rect 10968 14560 11020 14569
rect 4252 14424 4304 14433
rect 3976 14399 4028 14408
rect 3976 14365 3985 14399
rect 3985 14365 4019 14399
rect 4019 14365 4028 14399
rect 3976 14356 4028 14365
rect 4160 14399 4212 14408
rect 4160 14365 4169 14399
rect 4169 14365 4203 14399
rect 4203 14365 4212 14399
rect 4160 14356 4212 14365
rect 4528 14356 4580 14408
rect 3424 14288 3476 14340
rect 5172 14399 5224 14408
rect 5172 14365 5181 14399
rect 5181 14365 5215 14399
rect 5215 14365 5224 14399
rect 5172 14356 5224 14365
rect 5908 14399 5960 14408
rect 5908 14365 5917 14399
rect 5917 14365 5951 14399
rect 5951 14365 5960 14399
rect 5908 14356 5960 14365
rect 7196 14331 7248 14340
rect 3608 14220 3660 14272
rect 4988 14263 5040 14272
rect 4988 14229 4997 14263
rect 4997 14229 5031 14263
rect 5031 14229 5040 14263
rect 4988 14220 5040 14229
rect 5080 14220 5132 14272
rect 7196 14297 7205 14331
rect 7205 14297 7239 14331
rect 7239 14297 7248 14331
rect 7196 14288 7248 14297
rect 8024 14288 8076 14340
rect 8852 14424 8904 14476
rect 9220 14356 9272 14408
rect 12808 14603 12860 14612
rect 12808 14569 12817 14603
rect 12817 14569 12851 14603
rect 12851 14569 12860 14603
rect 12808 14560 12860 14569
rect 9680 14331 9732 14340
rect 9680 14297 9689 14331
rect 9689 14297 9723 14331
rect 9723 14297 9732 14331
rect 9680 14288 9732 14297
rect 6736 14220 6788 14272
rect 9772 14220 9824 14272
rect 10600 14331 10652 14340
rect 10600 14297 10609 14331
rect 10609 14297 10643 14331
rect 10643 14297 10652 14331
rect 10600 14288 10652 14297
rect 10784 14331 10836 14340
rect 10784 14297 10793 14331
rect 10793 14297 10827 14331
rect 10827 14297 10836 14331
rect 10784 14288 10836 14297
rect 10876 14288 10928 14340
rect 11060 14220 11112 14272
rect 12716 14220 12768 14272
rect 3519 14118 3571 14170
rect 3583 14118 3635 14170
rect 3647 14118 3699 14170
rect 3711 14118 3763 14170
rect 3775 14118 3827 14170
rect 7337 14118 7389 14170
rect 7401 14118 7453 14170
rect 7465 14118 7517 14170
rect 7529 14118 7581 14170
rect 7593 14118 7645 14170
rect 11155 14118 11207 14170
rect 11219 14118 11271 14170
rect 11283 14118 11335 14170
rect 11347 14118 11399 14170
rect 11411 14118 11463 14170
rect 14973 14118 15025 14170
rect 15037 14118 15089 14170
rect 15101 14118 15153 14170
rect 15165 14118 15217 14170
rect 15229 14118 15281 14170
rect 1400 13948 1452 14000
rect 1952 14016 2004 14068
rect 2228 14016 2280 14068
rect 2504 13948 2556 14000
rect 3240 14016 3292 14068
rect 3424 14016 3476 14068
rect 3976 14016 4028 14068
rect 5172 14016 5224 14068
rect 5908 14016 5960 14068
rect 6736 14059 6788 14068
rect 6736 14025 6745 14059
rect 6745 14025 6779 14059
rect 6779 14025 6788 14059
rect 6736 14016 6788 14025
rect 7288 14016 7340 14068
rect 7748 14016 7800 14068
rect 8944 14059 8996 14068
rect 8944 14025 8953 14059
rect 8953 14025 8987 14059
rect 8987 14025 8996 14059
rect 8944 14016 8996 14025
rect 1952 13855 2004 13864
rect 1952 13821 1961 13855
rect 1961 13821 1995 13855
rect 1995 13821 2004 13855
rect 1952 13812 2004 13821
rect 2228 13923 2280 13932
rect 2228 13889 2237 13923
rect 2237 13889 2271 13923
rect 2271 13889 2280 13923
rect 2228 13880 2280 13889
rect 7196 13948 7248 14000
rect 9220 13991 9272 14000
rect 2688 13812 2740 13864
rect 3424 13880 3476 13932
rect 4252 13880 4304 13932
rect 5080 13880 5132 13932
rect 2780 13744 2832 13796
rect 1860 13719 1912 13728
rect 1860 13685 1869 13719
rect 1869 13685 1903 13719
rect 1903 13685 1912 13719
rect 1860 13676 1912 13685
rect 1952 13676 2004 13728
rect 4160 13719 4212 13728
rect 4160 13685 4169 13719
rect 4169 13685 4203 13719
rect 4203 13685 4212 13719
rect 4160 13676 4212 13685
rect 4988 13812 5040 13864
rect 5356 13812 5408 13864
rect 7104 13923 7156 13932
rect 7104 13889 7113 13923
rect 7113 13889 7147 13923
rect 7147 13889 7156 13923
rect 7104 13880 7156 13889
rect 7564 13923 7616 13932
rect 7564 13889 7573 13923
rect 7573 13889 7607 13923
rect 7607 13889 7616 13923
rect 7564 13880 7616 13889
rect 7656 13923 7708 13932
rect 7656 13889 7665 13923
rect 7665 13889 7699 13923
rect 7699 13889 7708 13923
rect 7656 13880 7708 13889
rect 5264 13744 5316 13796
rect 6552 13744 6604 13796
rect 7196 13744 7248 13796
rect 8024 13812 8076 13864
rect 8392 13812 8444 13864
rect 8576 13812 8628 13864
rect 9220 13957 9229 13991
rect 9229 13957 9263 13991
rect 9263 13957 9272 13991
rect 9220 13948 9272 13957
rect 9128 13880 9180 13932
rect 8852 13812 8904 13864
rect 9680 14016 9732 14068
rect 9772 14016 9824 14068
rect 10876 14059 10928 14068
rect 10876 14025 10885 14059
rect 10885 14025 10919 14059
rect 10919 14025 10928 14059
rect 10876 14016 10928 14025
rect 10600 13880 10652 13932
rect 10876 13923 10928 13932
rect 10876 13889 10885 13923
rect 10885 13889 10919 13923
rect 10919 13889 10928 13923
rect 10876 13880 10928 13889
rect 6000 13676 6052 13728
rect 2859 13574 2911 13626
rect 2923 13574 2975 13626
rect 2987 13574 3039 13626
rect 3051 13574 3103 13626
rect 3115 13574 3167 13626
rect 6677 13574 6729 13626
rect 6741 13574 6793 13626
rect 6805 13574 6857 13626
rect 6869 13574 6921 13626
rect 6933 13574 6985 13626
rect 10495 13574 10547 13626
rect 10559 13574 10611 13626
rect 10623 13574 10675 13626
rect 10687 13574 10739 13626
rect 10751 13574 10803 13626
rect 14313 13574 14365 13626
rect 14377 13574 14429 13626
rect 14441 13574 14493 13626
rect 14505 13574 14557 13626
rect 14569 13574 14621 13626
rect 2596 13472 2648 13524
rect 2780 13472 2832 13524
rect 5264 13472 5316 13524
rect 5356 13472 5408 13524
rect 7012 13515 7064 13524
rect 7012 13481 7021 13515
rect 7021 13481 7055 13515
rect 7055 13481 7064 13515
rect 7012 13472 7064 13481
rect 7288 13472 7340 13524
rect 7564 13472 7616 13524
rect 8392 13515 8444 13524
rect 8392 13481 8401 13515
rect 8401 13481 8435 13515
rect 8435 13481 8444 13515
rect 8392 13472 8444 13481
rect 8576 13515 8628 13524
rect 8576 13481 8585 13515
rect 8585 13481 8619 13515
rect 8619 13481 8628 13515
rect 8576 13472 8628 13481
rect 9128 13472 9180 13524
rect 12348 13472 12400 13524
rect 12992 13472 13044 13524
rect 13912 13472 13964 13524
rect 1860 13336 1912 13388
rect 2136 13379 2188 13388
rect 2136 13345 2145 13379
rect 2145 13345 2179 13379
rect 2179 13345 2188 13379
rect 2136 13336 2188 13345
rect 940 13268 992 13320
rect 1952 13200 2004 13252
rect 2228 13311 2280 13320
rect 2228 13277 2237 13311
rect 2237 13277 2271 13311
rect 2271 13277 2280 13311
rect 2228 13268 2280 13277
rect 3240 13311 3292 13320
rect 3240 13277 3249 13311
rect 3249 13277 3283 13311
rect 3283 13277 3292 13311
rect 3240 13268 3292 13277
rect 2504 13200 2556 13252
rect 4160 13268 4212 13320
rect 5540 13268 5592 13320
rect 5908 13268 5960 13320
rect 7104 13404 7156 13456
rect 7380 13404 7432 13456
rect 7196 13268 7248 13320
rect 11060 13404 11112 13456
rect 2412 13175 2464 13184
rect 2412 13141 2421 13175
rect 2421 13141 2455 13175
rect 2455 13141 2464 13175
rect 2412 13132 2464 13141
rect 4896 13175 4948 13184
rect 4896 13141 4905 13175
rect 4905 13141 4939 13175
rect 4939 13141 4948 13175
rect 4896 13132 4948 13141
rect 6460 13132 6512 13184
rect 6552 13175 6604 13184
rect 6552 13141 6561 13175
rect 6561 13141 6595 13175
rect 6595 13141 6604 13175
rect 6552 13132 6604 13141
rect 7656 13311 7708 13320
rect 7656 13277 7665 13311
rect 7665 13277 7699 13311
rect 7699 13277 7708 13311
rect 7656 13268 7708 13277
rect 8392 13268 8444 13320
rect 10140 13311 10192 13320
rect 10140 13277 10149 13311
rect 10149 13277 10183 13311
rect 10183 13277 10192 13311
rect 10140 13268 10192 13277
rect 10692 13311 10744 13320
rect 10692 13277 10701 13311
rect 10701 13277 10735 13311
rect 10735 13277 10744 13311
rect 10692 13268 10744 13277
rect 10876 13311 10928 13320
rect 10876 13277 10885 13311
rect 10885 13277 10919 13311
rect 10919 13277 10928 13311
rect 10876 13268 10928 13277
rect 11520 13268 11572 13320
rect 11612 13311 11664 13320
rect 11612 13277 11621 13311
rect 11621 13277 11655 13311
rect 11655 13277 11664 13311
rect 11612 13268 11664 13277
rect 8300 13200 8352 13252
rect 8116 13132 8168 13184
rect 10324 13243 10376 13252
rect 10324 13209 10333 13243
rect 10333 13209 10367 13243
rect 10367 13209 10376 13243
rect 10324 13200 10376 13209
rect 12716 13311 12768 13320
rect 12716 13277 12725 13311
rect 12725 13277 12759 13311
rect 12759 13277 12768 13311
rect 12716 13268 12768 13277
rect 13912 13268 13964 13320
rect 15752 13311 15804 13320
rect 15752 13277 15761 13311
rect 15761 13277 15795 13311
rect 15795 13277 15804 13311
rect 15752 13268 15804 13277
rect 13636 13175 13688 13184
rect 13636 13141 13645 13175
rect 13645 13141 13679 13175
rect 13679 13141 13688 13175
rect 13636 13132 13688 13141
rect 14372 13132 14424 13184
rect 14832 13132 14884 13184
rect 15936 13175 15988 13184
rect 15936 13141 15945 13175
rect 15945 13141 15979 13175
rect 15979 13141 15988 13175
rect 15936 13132 15988 13141
rect 3519 13030 3571 13082
rect 3583 13030 3635 13082
rect 3647 13030 3699 13082
rect 3711 13030 3763 13082
rect 3775 13030 3827 13082
rect 7337 13030 7389 13082
rect 7401 13030 7453 13082
rect 7465 13030 7517 13082
rect 7529 13030 7581 13082
rect 7593 13030 7645 13082
rect 11155 13030 11207 13082
rect 11219 13030 11271 13082
rect 11283 13030 11335 13082
rect 11347 13030 11399 13082
rect 11411 13030 11463 13082
rect 14973 13030 15025 13082
rect 15037 13030 15089 13082
rect 15101 13030 15153 13082
rect 15165 13030 15217 13082
rect 15229 13030 15281 13082
rect 2504 12928 2556 12980
rect 2688 12971 2740 12980
rect 2688 12937 2697 12971
rect 2697 12937 2731 12971
rect 2731 12937 2740 12971
rect 2688 12928 2740 12937
rect 3240 12928 3292 12980
rect 4896 12928 4948 12980
rect 4988 12928 5040 12980
rect 5540 12971 5592 12980
rect 5540 12937 5549 12971
rect 5549 12937 5583 12971
rect 5583 12937 5592 12971
rect 5540 12928 5592 12937
rect 6552 12928 6604 12980
rect 8116 12928 8168 12980
rect 8300 12971 8352 12980
rect 8300 12937 8309 12971
rect 8309 12937 8343 12971
rect 8343 12937 8352 12971
rect 8300 12928 8352 12937
rect 8852 12928 8904 12980
rect 10140 12928 10192 12980
rect 10692 12928 10744 12980
rect 11520 12928 11572 12980
rect 15752 12928 15804 12980
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 5724 12835 5776 12844
rect 5724 12801 5733 12835
rect 5733 12801 5767 12835
rect 5767 12801 5776 12835
rect 5724 12792 5776 12801
rect 1860 12724 1912 12776
rect 2044 12724 2096 12776
rect 1676 12588 1728 12640
rect 2228 12588 2280 12640
rect 4252 12588 4304 12640
rect 6552 12588 6604 12640
rect 7104 12724 7156 12776
rect 7472 12792 7524 12844
rect 7288 12724 7340 12776
rect 7840 12792 7892 12844
rect 7932 12835 7984 12844
rect 7932 12801 7941 12835
rect 7941 12801 7975 12835
rect 7975 12801 7984 12835
rect 7932 12792 7984 12801
rect 9128 12860 9180 12912
rect 8300 12792 8352 12844
rect 10324 12835 10376 12844
rect 10324 12801 10333 12835
rect 10333 12801 10367 12835
rect 10367 12801 10376 12835
rect 10324 12792 10376 12801
rect 13636 12792 13688 12844
rect 14832 12792 14884 12844
rect 8300 12656 8352 12708
rect 10048 12724 10100 12776
rect 11612 12767 11664 12776
rect 11612 12733 11621 12767
rect 11621 12733 11655 12767
rect 11655 12733 11664 12767
rect 11612 12724 11664 12733
rect 13360 12767 13412 12776
rect 13360 12733 13369 12767
rect 13369 12733 13403 12767
rect 13403 12733 13412 12767
rect 13360 12724 13412 12733
rect 14372 12724 14424 12776
rect 7840 12588 7892 12640
rect 8576 12631 8628 12640
rect 8576 12597 8585 12631
rect 8585 12597 8619 12631
rect 8619 12597 8628 12631
rect 8576 12588 8628 12597
rect 12072 12631 12124 12640
rect 12072 12597 12081 12631
rect 12081 12597 12115 12631
rect 12115 12597 12124 12631
rect 12072 12588 12124 12597
rect 2859 12486 2911 12538
rect 2923 12486 2975 12538
rect 2987 12486 3039 12538
rect 3051 12486 3103 12538
rect 3115 12486 3167 12538
rect 6677 12486 6729 12538
rect 6741 12486 6793 12538
rect 6805 12486 6857 12538
rect 6869 12486 6921 12538
rect 6933 12486 6985 12538
rect 10495 12486 10547 12538
rect 10559 12486 10611 12538
rect 10623 12486 10675 12538
rect 10687 12486 10739 12538
rect 10751 12486 10803 12538
rect 14313 12486 14365 12538
rect 14377 12486 14429 12538
rect 14441 12486 14493 12538
rect 14505 12486 14557 12538
rect 14569 12486 14621 12538
rect 2044 12427 2096 12436
rect 2044 12393 2053 12427
rect 2053 12393 2087 12427
rect 2087 12393 2096 12427
rect 2044 12384 2096 12393
rect 5080 12384 5132 12436
rect 5724 12384 5776 12436
rect 5908 12427 5960 12436
rect 5908 12393 5917 12427
rect 5917 12393 5951 12427
rect 5951 12393 5960 12427
rect 5908 12384 5960 12393
rect 8392 12384 8444 12436
rect 10048 12384 10100 12436
rect 12348 12427 12400 12436
rect 12348 12393 12357 12427
rect 12357 12393 12391 12427
rect 12391 12393 12400 12427
rect 12348 12384 12400 12393
rect 1676 12223 1728 12232
rect 1676 12189 1685 12223
rect 1685 12189 1719 12223
rect 1719 12189 1728 12223
rect 1676 12180 1728 12189
rect 2504 12223 2556 12232
rect 2504 12189 2513 12223
rect 2513 12189 2547 12223
rect 2547 12189 2556 12223
rect 2504 12180 2556 12189
rect 3424 12223 3476 12232
rect 3424 12189 3433 12223
rect 3433 12189 3467 12223
rect 3467 12189 3476 12223
rect 3424 12180 3476 12189
rect 4160 12180 4212 12232
rect 4252 12223 4304 12232
rect 4252 12189 4261 12223
rect 4261 12189 4295 12223
rect 4295 12189 4304 12223
rect 4252 12180 4304 12189
rect 4712 12223 4764 12232
rect 4712 12189 4721 12223
rect 4721 12189 4755 12223
rect 4755 12189 4764 12223
rect 4712 12180 4764 12189
rect 1952 12112 2004 12164
rect 2228 12112 2280 12164
rect 3240 12155 3292 12164
rect 3240 12121 3249 12155
rect 3249 12121 3283 12155
rect 3283 12121 3292 12155
rect 5908 12223 5960 12232
rect 5908 12189 5917 12223
rect 5917 12189 5951 12223
rect 5951 12189 5960 12223
rect 5908 12180 5960 12189
rect 6000 12180 6052 12232
rect 6184 12223 6236 12232
rect 6184 12189 6193 12223
rect 6193 12189 6227 12223
rect 6227 12189 6236 12223
rect 6184 12180 6236 12189
rect 7104 12316 7156 12368
rect 8024 12316 8076 12368
rect 11980 12359 12032 12368
rect 11980 12325 11989 12359
rect 11989 12325 12023 12359
rect 12023 12325 12032 12359
rect 11980 12316 12032 12325
rect 7748 12248 7800 12300
rect 9036 12291 9088 12300
rect 9036 12257 9045 12291
rect 9045 12257 9079 12291
rect 9079 12257 9088 12291
rect 9036 12248 9088 12257
rect 7472 12180 7524 12232
rect 7840 12223 7892 12232
rect 7840 12189 7849 12223
rect 7849 12189 7883 12223
rect 7883 12189 7892 12223
rect 7840 12180 7892 12189
rect 3240 12112 3292 12121
rect 6552 12112 6604 12164
rect 8024 12223 8076 12232
rect 8024 12189 8033 12223
rect 8033 12189 8067 12223
rect 8067 12189 8076 12223
rect 8024 12180 8076 12189
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 12072 12180 12124 12232
rect 13912 12427 13964 12436
rect 13912 12393 13921 12427
rect 13921 12393 13955 12427
rect 13955 12393 13964 12427
rect 13912 12384 13964 12393
rect 13636 12316 13688 12368
rect 4068 12087 4120 12096
rect 4068 12053 4077 12087
rect 4077 12053 4111 12087
rect 4111 12053 4120 12087
rect 4068 12044 4120 12053
rect 9956 12044 10008 12096
rect 10876 12044 10928 12096
rect 13452 12155 13504 12164
rect 13452 12121 13461 12155
rect 13461 12121 13495 12155
rect 13495 12121 13504 12155
rect 13452 12112 13504 12121
rect 12900 12087 12952 12096
rect 12900 12053 12909 12087
rect 12909 12053 12943 12087
rect 12943 12053 12952 12087
rect 12900 12044 12952 12053
rect 3519 11942 3571 11994
rect 3583 11942 3635 11994
rect 3647 11942 3699 11994
rect 3711 11942 3763 11994
rect 3775 11942 3827 11994
rect 7337 11942 7389 11994
rect 7401 11942 7453 11994
rect 7465 11942 7517 11994
rect 7529 11942 7581 11994
rect 7593 11942 7645 11994
rect 11155 11942 11207 11994
rect 11219 11942 11271 11994
rect 11283 11942 11335 11994
rect 11347 11942 11399 11994
rect 11411 11942 11463 11994
rect 14973 11942 15025 11994
rect 15037 11942 15089 11994
rect 15101 11942 15153 11994
rect 15165 11942 15217 11994
rect 15229 11942 15281 11994
rect 3240 11840 3292 11892
rect 3424 11840 3476 11892
rect 4068 11840 4120 11892
rect 4712 11840 4764 11892
rect 4252 11772 4304 11824
rect 7196 11772 7248 11824
rect 7564 11772 7616 11824
rect 4160 11747 4212 11756
rect 4160 11713 4169 11747
rect 4169 11713 4203 11747
rect 4203 11713 4212 11747
rect 4160 11704 4212 11713
rect 9036 11840 9088 11892
rect 8852 11772 8904 11824
rect 8484 11636 8536 11688
rect 3884 11543 3936 11552
rect 3884 11509 3893 11543
rect 3893 11509 3927 11543
rect 3927 11509 3936 11543
rect 3884 11500 3936 11509
rect 6644 11500 6696 11552
rect 7472 11500 7524 11552
rect 7656 11500 7708 11552
rect 8576 11543 8628 11552
rect 8576 11509 8585 11543
rect 8585 11509 8619 11543
rect 8619 11509 8628 11543
rect 8576 11500 8628 11509
rect 8668 11500 8720 11552
rect 9956 11704 10008 11756
rect 10876 11883 10928 11892
rect 10876 11849 10885 11883
rect 10885 11849 10919 11883
rect 10919 11849 10928 11883
rect 10876 11840 10928 11849
rect 11980 11840 12032 11892
rect 12256 11840 12308 11892
rect 12900 11840 12952 11892
rect 14832 11883 14884 11892
rect 14832 11849 14841 11883
rect 14841 11849 14875 11883
rect 14875 11849 14884 11883
rect 14832 11840 14884 11849
rect 9680 11568 9732 11620
rect 11520 11747 11572 11756
rect 11520 11713 11529 11747
rect 11529 11713 11563 11747
rect 11563 11713 11572 11747
rect 11520 11704 11572 11713
rect 11704 11747 11756 11756
rect 11704 11713 11713 11747
rect 11713 11713 11747 11747
rect 11747 11713 11756 11747
rect 11704 11704 11756 11713
rect 14096 11704 14148 11756
rect 14832 11704 14884 11756
rect 15016 11747 15068 11756
rect 15016 11713 15025 11747
rect 15025 11713 15059 11747
rect 15059 11713 15068 11747
rect 15016 11704 15068 11713
rect 15200 11636 15252 11688
rect 14188 11500 14240 11552
rect 2859 11398 2911 11450
rect 2923 11398 2975 11450
rect 2987 11398 3039 11450
rect 3051 11398 3103 11450
rect 3115 11398 3167 11450
rect 6677 11398 6729 11450
rect 6741 11398 6793 11450
rect 6805 11398 6857 11450
rect 6869 11398 6921 11450
rect 6933 11398 6985 11450
rect 10495 11398 10547 11450
rect 10559 11398 10611 11450
rect 10623 11398 10675 11450
rect 10687 11398 10739 11450
rect 10751 11398 10803 11450
rect 14313 11398 14365 11450
rect 14377 11398 14429 11450
rect 14441 11398 14493 11450
rect 14505 11398 14557 11450
rect 14569 11398 14621 11450
rect 6460 11339 6512 11348
rect 6460 11305 6469 11339
rect 6469 11305 6503 11339
rect 6503 11305 6512 11339
rect 6460 11296 6512 11305
rect 7104 11296 7156 11348
rect 8668 11339 8720 11348
rect 8668 11305 8677 11339
rect 8677 11305 8711 11339
rect 8711 11305 8720 11339
rect 8668 11296 8720 11305
rect 5816 11228 5868 11280
rect 6736 11160 6788 11212
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 7748 11228 7800 11280
rect 9680 11228 9732 11280
rect 11704 11228 11756 11280
rect 7104 11067 7156 11076
rect 7104 11033 7113 11067
rect 7113 11033 7147 11067
rect 7147 11033 7156 11067
rect 7104 11024 7156 11033
rect 7472 11135 7524 11144
rect 7472 11101 7481 11135
rect 7481 11101 7515 11135
rect 7515 11101 7524 11135
rect 7472 11092 7524 11101
rect 7564 11135 7616 11144
rect 7564 11101 7573 11135
rect 7573 11101 7607 11135
rect 7607 11101 7616 11135
rect 7564 11092 7616 11101
rect 7656 11092 7708 11144
rect 8484 11092 8536 11144
rect 8852 11092 8904 11144
rect 7748 11067 7800 11076
rect 7748 11033 7757 11067
rect 7757 11033 7791 11067
rect 7791 11033 7800 11067
rect 7748 11024 7800 11033
rect 11520 11092 11572 11144
rect 15016 11296 15068 11348
rect 15200 11296 15252 11348
rect 12256 11092 12308 11144
rect 13820 11228 13872 11280
rect 13544 11160 13596 11212
rect 14188 11160 14240 11212
rect 13360 11135 13412 11144
rect 13360 11101 13369 11135
rect 13369 11101 13403 11135
rect 13403 11101 13412 11135
rect 13360 11092 13412 11101
rect 14096 11092 14148 11144
rect 15660 11203 15712 11212
rect 15660 11169 15669 11203
rect 15669 11169 15703 11203
rect 15703 11169 15712 11203
rect 15660 11160 15712 11169
rect 14832 11092 14884 11144
rect 6184 10956 6236 11008
rect 6276 10956 6328 11008
rect 6460 10956 6512 11008
rect 7472 10956 7524 11008
rect 7932 10956 7984 11008
rect 9680 10956 9732 11008
rect 14004 11024 14056 11076
rect 3519 10854 3571 10906
rect 3583 10854 3635 10906
rect 3647 10854 3699 10906
rect 3711 10854 3763 10906
rect 3775 10854 3827 10906
rect 7337 10854 7389 10906
rect 7401 10854 7453 10906
rect 7465 10854 7517 10906
rect 7529 10854 7581 10906
rect 7593 10854 7645 10906
rect 11155 10854 11207 10906
rect 11219 10854 11271 10906
rect 11283 10854 11335 10906
rect 11347 10854 11399 10906
rect 11411 10854 11463 10906
rect 14973 10854 15025 10906
rect 15037 10854 15089 10906
rect 15101 10854 15153 10906
rect 15165 10854 15217 10906
rect 15229 10854 15281 10906
rect 3884 10752 3936 10804
rect 4160 10752 4212 10804
rect 2412 10684 2464 10736
rect 5724 10752 5776 10804
rect 6092 10752 6144 10804
rect 9956 10752 10008 10804
rect 13452 10752 13504 10804
rect 16028 10752 16080 10804
rect 940 10616 992 10668
rect 4620 10684 4672 10736
rect 6368 10684 6420 10736
rect 2412 10591 2464 10600
rect 2412 10557 2421 10591
rect 2421 10557 2455 10591
rect 2455 10557 2464 10591
rect 2412 10548 2464 10557
rect 4436 10480 4488 10532
rect 5080 10616 5132 10668
rect 3424 10412 3476 10464
rect 3608 10412 3660 10464
rect 3884 10455 3936 10464
rect 3884 10421 3893 10455
rect 3893 10421 3927 10455
rect 3927 10421 3936 10455
rect 3884 10412 3936 10421
rect 4344 10412 4396 10464
rect 5632 10412 5684 10464
rect 6000 10659 6052 10668
rect 6000 10625 6009 10659
rect 6009 10625 6043 10659
rect 6043 10625 6052 10659
rect 6000 10616 6052 10625
rect 6092 10659 6144 10668
rect 6092 10625 6101 10659
rect 6101 10625 6135 10659
rect 6135 10625 6144 10659
rect 6092 10616 6144 10625
rect 6552 10616 6604 10668
rect 5908 10591 5960 10600
rect 5908 10557 5917 10591
rect 5917 10557 5951 10591
rect 5951 10557 5960 10591
rect 5908 10548 5960 10557
rect 6276 10548 6328 10600
rect 7104 10548 7156 10600
rect 12348 10548 12400 10600
rect 12716 10659 12768 10668
rect 12716 10625 12725 10659
rect 12725 10625 12759 10659
rect 12759 10625 12768 10659
rect 12716 10616 12768 10625
rect 13544 10684 13596 10736
rect 15660 10727 15712 10736
rect 15660 10693 15669 10727
rect 15669 10693 15703 10727
rect 15703 10693 15712 10727
rect 15660 10684 15712 10693
rect 13360 10548 13412 10600
rect 7748 10412 7800 10464
rect 8300 10412 8352 10464
rect 8392 10412 8444 10464
rect 9312 10412 9364 10464
rect 2859 10310 2911 10362
rect 2923 10310 2975 10362
rect 2987 10310 3039 10362
rect 3051 10310 3103 10362
rect 3115 10310 3167 10362
rect 6677 10310 6729 10362
rect 6741 10310 6793 10362
rect 6805 10310 6857 10362
rect 6869 10310 6921 10362
rect 6933 10310 6985 10362
rect 10495 10310 10547 10362
rect 10559 10310 10611 10362
rect 10623 10310 10675 10362
rect 10687 10310 10739 10362
rect 10751 10310 10803 10362
rect 14313 10310 14365 10362
rect 14377 10310 14429 10362
rect 14441 10310 14493 10362
rect 14505 10310 14557 10362
rect 14569 10310 14621 10362
rect 2412 10208 2464 10260
rect 3884 10208 3936 10260
rect 3608 10140 3660 10192
rect 5540 10208 5592 10260
rect 6000 10251 6052 10260
rect 6000 10217 6009 10251
rect 6009 10217 6043 10251
rect 6043 10217 6052 10251
rect 6000 10208 6052 10217
rect 6092 10208 6144 10260
rect 8392 10208 8444 10260
rect 9496 10208 9548 10260
rect 4344 10140 4396 10192
rect 1492 9911 1544 9920
rect 1492 9877 1501 9911
rect 1501 9877 1535 9911
rect 1535 9877 1544 9911
rect 1492 9868 1544 9877
rect 3240 10047 3292 10056
rect 3240 10013 3249 10047
rect 3249 10013 3283 10047
rect 3283 10013 3292 10047
rect 3240 10004 3292 10013
rect 4436 10047 4488 10056
rect 4436 10013 4445 10047
rect 4445 10013 4479 10047
rect 4479 10013 4488 10047
rect 4436 10004 4488 10013
rect 4620 10004 4672 10056
rect 5908 10140 5960 10192
rect 9680 10140 9732 10192
rect 9956 10140 10008 10192
rect 5080 10047 5132 10056
rect 5080 10013 5089 10047
rect 5089 10013 5123 10047
rect 5123 10013 5132 10047
rect 5080 10004 5132 10013
rect 5632 10072 5684 10124
rect 5724 10004 5776 10056
rect 5816 10004 5868 10056
rect 6368 10072 6420 10124
rect 6092 10047 6144 10056
rect 6092 10013 6101 10047
rect 6101 10013 6135 10047
rect 6135 10013 6144 10047
rect 6092 10004 6144 10013
rect 6460 10004 6512 10056
rect 6552 10047 6604 10056
rect 6552 10013 6561 10047
rect 6561 10013 6595 10047
rect 6595 10013 6604 10047
rect 6552 10004 6604 10013
rect 12348 10251 12400 10260
rect 12348 10217 12357 10251
rect 12357 10217 12391 10251
rect 12391 10217 12400 10251
rect 12348 10208 12400 10217
rect 12716 10251 12768 10260
rect 12716 10217 12725 10251
rect 12725 10217 12759 10251
rect 12759 10217 12768 10251
rect 12716 10208 12768 10217
rect 14832 10208 14884 10260
rect 6920 10047 6972 10056
rect 6920 10013 6929 10047
rect 6929 10013 6963 10047
rect 6963 10013 6972 10047
rect 6920 10004 6972 10013
rect 9036 10004 9088 10056
rect 9312 10047 9364 10056
rect 9312 10013 9321 10047
rect 9321 10013 9355 10047
rect 9355 10013 9364 10047
rect 9312 10004 9364 10013
rect 4160 9868 4212 9920
rect 5908 9868 5960 9920
rect 8116 9979 8168 9988
rect 8116 9945 8125 9979
rect 8125 9945 8159 9979
rect 8159 9945 8168 9979
rect 8116 9936 8168 9945
rect 8576 9936 8628 9988
rect 8208 9868 8260 9920
rect 9496 10004 9548 10056
rect 9956 10004 10008 10056
rect 10324 9936 10376 9988
rect 12072 10004 12124 10056
rect 14832 10004 14884 10056
rect 11520 9868 11572 9920
rect 12256 9868 12308 9920
rect 15660 9979 15712 9988
rect 15660 9945 15669 9979
rect 15669 9945 15703 9979
rect 15703 9945 15712 9979
rect 15660 9936 15712 9945
rect 15384 9868 15436 9920
rect 15568 9868 15620 9920
rect 16028 9868 16080 9920
rect 3519 9766 3571 9818
rect 3583 9766 3635 9818
rect 3647 9766 3699 9818
rect 3711 9766 3763 9818
rect 3775 9766 3827 9818
rect 7337 9766 7389 9818
rect 7401 9766 7453 9818
rect 7465 9766 7517 9818
rect 7529 9766 7581 9818
rect 7593 9766 7645 9818
rect 11155 9766 11207 9818
rect 11219 9766 11271 9818
rect 11283 9766 11335 9818
rect 11347 9766 11399 9818
rect 11411 9766 11463 9818
rect 14973 9766 15025 9818
rect 15037 9766 15089 9818
rect 15101 9766 15153 9818
rect 15165 9766 15217 9818
rect 15229 9766 15281 9818
rect 3240 9664 3292 9716
rect 3424 9664 3476 9716
rect 7012 9664 7064 9716
rect 1676 9528 1728 9580
rect 4344 9639 4396 9648
rect 3332 9528 3384 9580
rect 4344 9605 4353 9639
rect 4353 9605 4387 9639
rect 4387 9605 4396 9639
rect 4344 9596 4396 9605
rect 4528 9596 4580 9648
rect 6920 9596 6972 9648
rect 7564 9596 7616 9648
rect 8208 9664 8260 9716
rect 8116 9596 8168 9648
rect 8392 9596 8444 9648
rect 8576 9596 8628 9648
rect 9036 9639 9088 9648
rect 9036 9605 9045 9639
rect 9045 9605 9079 9639
rect 9079 9605 9088 9639
rect 9036 9596 9088 9605
rect 7196 9460 7248 9512
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 7656 9528 7708 9580
rect 7472 9392 7524 9444
rect 3884 9367 3936 9376
rect 3884 9333 3893 9367
rect 3893 9333 3927 9367
rect 3927 9333 3936 9367
rect 3884 9324 3936 9333
rect 6460 9324 6512 9376
rect 9128 9528 9180 9580
rect 10324 9528 10376 9580
rect 13360 9707 13412 9716
rect 13360 9673 13369 9707
rect 13369 9673 13403 9707
rect 13403 9673 13412 9707
rect 13360 9664 13412 9673
rect 13912 9664 13964 9716
rect 13176 9571 13228 9580
rect 13176 9537 13185 9571
rect 13185 9537 13219 9571
rect 13219 9537 13228 9571
rect 13176 9528 13228 9537
rect 13636 9528 13688 9580
rect 14004 9528 14056 9580
rect 14648 9528 14700 9580
rect 15384 9528 15436 9580
rect 9956 9392 10008 9444
rect 10508 9503 10560 9512
rect 10508 9469 10517 9503
rect 10517 9469 10551 9503
rect 10551 9469 10560 9503
rect 10508 9460 10560 9469
rect 11520 9503 11572 9512
rect 8024 9324 8076 9376
rect 9312 9324 9364 9376
rect 10324 9324 10376 9376
rect 11520 9469 11529 9503
rect 11529 9469 11563 9503
rect 11563 9469 11572 9503
rect 11520 9460 11572 9469
rect 14740 9503 14792 9512
rect 14740 9469 14749 9503
rect 14749 9469 14783 9503
rect 14783 9469 14792 9503
rect 14740 9460 14792 9469
rect 15568 9503 15620 9512
rect 15568 9469 15577 9503
rect 15577 9469 15611 9503
rect 15611 9469 15620 9503
rect 15568 9460 15620 9469
rect 15660 9460 15712 9512
rect 11888 9367 11940 9376
rect 11888 9333 11897 9367
rect 11897 9333 11931 9367
rect 11931 9333 11940 9367
rect 11888 9324 11940 9333
rect 2859 9222 2911 9274
rect 2923 9222 2975 9274
rect 2987 9222 3039 9274
rect 3051 9222 3103 9274
rect 3115 9222 3167 9274
rect 6677 9222 6729 9274
rect 6741 9222 6793 9274
rect 6805 9222 6857 9274
rect 6869 9222 6921 9274
rect 6933 9222 6985 9274
rect 10495 9222 10547 9274
rect 10559 9222 10611 9274
rect 10623 9222 10675 9274
rect 10687 9222 10739 9274
rect 10751 9222 10803 9274
rect 14313 9222 14365 9274
rect 14377 9222 14429 9274
rect 14441 9222 14493 9274
rect 14505 9222 14557 9274
rect 14569 9222 14621 9274
rect 4344 9120 4396 9172
rect 9772 9120 9824 9172
rect 11888 9120 11940 9172
rect 12256 9120 12308 9172
rect 13176 9163 13228 9172
rect 13176 9129 13185 9163
rect 13185 9129 13219 9163
rect 13219 9129 13228 9163
rect 13176 9120 13228 9129
rect 14740 9120 14792 9172
rect 14832 9163 14884 9172
rect 14832 9129 14841 9163
rect 14841 9129 14875 9163
rect 14875 9129 14884 9163
rect 14832 9120 14884 9129
rect 5908 9052 5960 9104
rect 6184 8984 6236 9036
rect 5540 8916 5592 8968
rect 6552 9052 6604 9104
rect 7472 9095 7524 9104
rect 7472 9061 7481 9095
rect 7481 9061 7515 9095
rect 7515 9061 7524 9095
rect 7472 9052 7524 9061
rect 6552 8959 6604 8968
rect 6552 8925 6561 8959
rect 6561 8925 6595 8959
rect 6595 8925 6604 8959
rect 6552 8916 6604 8925
rect 6736 8959 6788 8968
rect 6736 8925 6745 8959
rect 6745 8925 6779 8959
rect 6779 8925 6788 8959
rect 6736 8916 6788 8925
rect 7656 8984 7708 9036
rect 8116 9027 8168 9036
rect 8116 8993 8125 9027
rect 8125 8993 8159 9027
rect 8159 8993 8168 9027
rect 8116 8984 8168 8993
rect 8392 9052 8444 9104
rect 9128 9052 9180 9104
rect 7564 8959 7616 8968
rect 7564 8925 7573 8959
rect 7573 8925 7607 8959
rect 7607 8925 7616 8959
rect 7564 8916 7616 8925
rect 940 8848 992 8900
rect 1768 8891 1820 8900
rect 1768 8857 1777 8891
rect 1777 8857 1811 8891
rect 1811 8857 1820 8891
rect 1768 8848 1820 8857
rect 5724 8848 5776 8900
rect 6000 8848 6052 8900
rect 7840 8780 7892 8832
rect 8392 8916 8444 8968
rect 8576 8916 8628 8968
rect 12164 9095 12216 9104
rect 12164 9061 12173 9095
rect 12173 9061 12207 9095
rect 12207 9061 12216 9095
rect 12164 9052 12216 9061
rect 11520 8916 11572 8968
rect 8300 8780 8352 8832
rect 12164 8848 12216 8900
rect 14648 8959 14700 8968
rect 14648 8925 14657 8959
rect 14657 8925 14691 8959
rect 14691 8925 14700 8959
rect 14648 8916 14700 8925
rect 11704 8780 11756 8832
rect 3519 8678 3571 8730
rect 3583 8678 3635 8730
rect 3647 8678 3699 8730
rect 3711 8678 3763 8730
rect 3775 8678 3827 8730
rect 7337 8678 7389 8730
rect 7401 8678 7453 8730
rect 7465 8678 7517 8730
rect 7529 8678 7581 8730
rect 7593 8678 7645 8730
rect 11155 8678 11207 8730
rect 11219 8678 11271 8730
rect 11283 8678 11335 8730
rect 11347 8678 11399 8730
rect 11411 8678 11463 8730
rect 14973 8678 15025 8730
rect 15037 8678 15089 8730
rect 15101 8678 15153 8730
rect 15165 8678 15217 8730
rect 15229 8678 15281 8730
rect 3516 8576 3568 8628
rect 3884 8576 3936 8628
rect 5540 8576 5592 8628
rect 6736 8576 6788 8628
rect 7748 8619 7800 8628
rect 7748 8585 7757 8619
rect 7757 8585 7791 8619
rect 7791 8585 7800 8619
rect 7748 8576 7800 8585
rect 8024 8576 8076 8628
rect 9036 8576 9088 8628
rect 10416 8576 10468 8628
rect 11520 8576 11572 8628
rect 12164 8576 12216 8628
rect 15384 8619 15436 8628
rect 15384 8585 15393 8619
rect 15393 8585 15427 8619
rect 15427 8585 15436 8619
rect 15384 8576 15436 8585
rect 2136 8483 2188 8492
rect 2136 8449 2145 8483
rect 2145 8449 2179 8483
rect 2179 8449 2188 8483
rect 2136 8440 2188 8449
rect 2596 8440 2648 8492
rect 3424 8483 3476 8492
rect 3424 8449 3433 8483
rect 3433 8449 3467 8483
rect 3467 8449 3476 8483
rect 3424 8440 3476 8449
rect 1952 8372 2004 8424
rect 2044 8372 2096 8424
rect 3884 8483 3936 8492
rect 3884 8449 3893 8483
rect 3893 8449 3927 8483
rect 3927 8449 3936 8483
rect 3884 8440 3936 8449
rect 4068 8440 4120 8492
rect 5540 8440 5592 8492
rect 5724 8483 5776 8492
rect 5724 8449 5733 8483
rect 5733 8449 5767 8483
rect 5767 8449 5776 8483
rect 5724 8440 5776 8449
rect 5908 8483 5960 8492
rect 5908 8449 5917 8483
rect 5917 8449 5951 8483
rect 5951 8449 5960 8483
rect 5908 8440 5960 8449
rect 6000 8483 6052 8492
rect 6000 8449 6009 8483
rect 6009 8449 6043 8483
rect 6043 8449 6052 8483
rect 6000 8440 6052 8449
rect 6552 8508 6604 8560
rect 6184 8483 6236 8492
rect 6184 8449 6193 8483
rect 6193 8449 6227 8483
rect 6227 8449 6236 8483
rect 8208 8508 8260 8560
rect 9312 8508 9364 8560
rect 6184 8440 6236 8449
rect 7472 8440 7524 8492
rect 2780 8347 2832 8356
rect 2780 8313 2789 8347
rect 2789 8313 2823 8347
rect 2823 8313 2832 8347
rect 2780 8304 2832 8313
rect 4436 8304 4488 8356
rect 2412 8236 2464 8288
rect 4252 8236 4304 8288
rect 7012 8372 7064 8424
rect 7288 8372 7340 8424
rect 10048 8483 10100 8492
rect 10048 8449 10057 8483
rect 10057 8449 10091 8483
rect 10091 8449 10100 8483
rect 10048 8440 10100 8449
rect 8944 8372 8996 8424
rect 9220 8372 9272 8424
rect 9680 8415 9732 8424
rect 9680 8381 9689 8415
rect 9689 8381 9723 8415
rect 9723 8381 9732 8415
rect 9680 8372 9732 8381
rect 11704 8483 11756 8492
rect 11704 8449 11713 8483
rect 11713 8449 11747 8483
rect 11747 8449 11756 8483
rect 11704 8440 11756 8449
rect 14740 8440 14792 8492
rect 14924 8483 14976 8492
rect 14924 8449 14933 8483
rect 14933 8449 14967 8483
rect 14967 8449 14976 8483
rect 14924 8440 14976 8449
rect 5632 8347 5684 8356
rect 5632 8313 5641 8347
rect 5641 8313 5675 8347
rect 5675 8313 5684 8347
rect 5632 8304 5684 8313
rect 7196 8304 7248 8356
rect 7012 8236 7064 8288
rect 14832 8372 14884 8424
rect 12440 8279 12492 8288
rect 12440 8245 12449 8279
rect 12449 8245 12483 8279
rect 12483 8245 12492 8279
rect 12440 8236 12492 8245
rect 2859 8134 2911 8186
rect 2923 8134 2975 8186
rect 2987 8134 3039 8186
rect 3051 8134 3103 8186
rect 3115 8134 3167 8186
rect 6677 8134 6729 8186
rect 6741 8134 6793 8186
rect 6805 8134 6857 8186
rect 6869 8134 6921 8186
rect 6933 8134 6985 8186
rect 10495 8134 10547 8186
rect 10559 8134 10611 8186
rect 10623 8134 10675 8186
rect 10687 8134 10739 8186
rect 10751 8134 10803 8186
rect 14313 8134 14365 8186
rect 14377 8134 14429 8186
rect 14441 8134 14493 8186
rect 14505 8134 14557 8186
rect 14569 8134 14621 8186
rect 1768 8032 1820 8084
rect 1952 8032 2004 8084
rect 2044 7964 2096 8016
rect 2596 8032 2648 8084
rect 2228 7964 2280 8016
rect 4620 8075 4672 8084
rect 4620 8041 4629 8075
rect 4629 8041 4663 8075
rect 4663 8041 4672 8075
rect 4620 8032 4672 8041
rect 5356 8032 5408 8084
rect 7840 8032 7892 8084
rect 8116 8032 8168 8084
rect 8392 8075 8444 8084
rect 8392 8041 8401 8075
rect 8401 8041 8435 8075
rect 8435 8041 8444 8075
rect 8392 8032 8444 8041
rect 8760 8032 8812 8084
rect 12256 8032 12308 8084
rect 5540 7964 5592 8016
rect 8944 7964 8996 8016
rect 9588 7964 9640 8016
rect 14924 8032 14976 8084
rect 1768 7692 1820 7744
rect 2228 7871 2280 7880
rect 2228 7837 2237 7871
rect 2237 7837 2271 7871
rect 2271 7837 2280 7871
rect 2228 7828 2280 7837
rect 2412 7896 2464 7948
rect 3424 7896 3476 7948
rect 3608 7896 3660 7948
rect 2596 7828 2648 7880
rect 2044 7803 2096 7812
rect 2044 7769 2061 7803
rect 2061 7769 2096 7803
rect 2044 7760 2096 7769
rect 3332 7828 3384 7880
rect 4620 7896 4672 7948
rect 9036 7939 9088 7948
rect 9036 7905 9045 7939
rect 9045 7905 9079 7939
rect 9079 7905 9088 7939
rect 9036 7896 9088 7905
rect 4344 7828 4396 7880
rect 4252 7760 4304 7812
rect 4896 7871 4948 7880
rect 4896 7837 4905 7871
rect 4905 7837 4939 7871
rect 4939 7837 4948 7871
rect 4896 7828 4948 7837
rect 6828 7871 6880 7880
rect 6828 7837 6837 7871
rect 6837 7837 6871 7871
rect 6871 7837 6880 7871
rect 6828 7828 6880 7837
rect 7012 7828 7064 7880
rect 7196 7828 7248 7880
rect 7472 7871 7524 7880
rect 7472 7837 7481 7871
rect 7481 7837 7515 7871
rect 7515 7837 7524 7871
rect 7472 7828 7524 7837
rect 2596 7692 2648 7744
rect 2872 7735 2924 7744
rect 2872 7701 2881 7735
rect 2881 7701 2915 7735
rect 2915 7701 2924 7735
rect 2872 7692 2924 7701
rect 3608 7692 3660 7744
rect 3976 7735 4028 7744
rect 3976 7701 3985 7735
rect 3985 7701 4019 7735
rect 4019 7701 4028 7735
rect 3976 7692 4028 7701
rect 4344 7692 4396 7744
rect 7288 7803 7340 7812
rect 7288 7769 7297 7803
rect 7297 7769 7331 7803
rect 7331 7769 7340 7803
rect 7288 7760 7340 7769
rect 8944 7871 8996 7880
rect 8944 7837 8953 7871
rect 8953 7837 8987 7871
rect 8987 7837 8996 7871
rect 8944 7828 8996 7837
rect 9312 7896 9364 7948
rect 9680 7939 9732 7948
rect 9680 7905 9689 7939
rect 9689 7905 9723 7939
rect 9723 7905 9732 7939
rect 9680 7896 9732 7905
rect 8024 7692 8076 7744
rect 8392 7692 8444 7744
rect 8576 7735 8628 7744
rect 8576 7701 8603 7735
rect 8603 7701 8628 7735
rect 8576 7692 8628 7701
rect 8668 7692 8720 7744
rect 9128 7760 9180 7812
rect 12072 7871 12124 7880
rect 12072 7837 12081 7871
rect 12081 7837 12115 7871
rect 12115 7837 12124 7871
rect 12072 7828 12124 7837
rect 12440 7828 12492 7880
rect 13176 7896 13228 7948
rect 14372 7939 14424 7948
rect 14372 7905 14381 7939
rect 14381 7905 14415 7939
rect 14415 7905 14424 7939
rect 14372 7896 14424 7905
rect 12900 7871 12952 7880
rect 12900 7837 12909 7871
rect 12909 7837 12943 7871
rect 12943 7837 12952 7871
rect 12900 7828 12952 7837
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 13820 7828 13872 7880
rect 14464 7871 14516 7880
rect 14464 7837 14473 7871
rect 14473 7837 14507 7871
rect 14507 7837 14516 7871
rect 14464 7828 14516 7837
rect 14740 7828 14792 7880
rect 12164 7735 12216 7744
rect 12164 7701 12173 7735
rect 12173 7701 12207 7735
rect 12207 7701 12216 7735
rect 12164 7692 12216 7701
rect 15936 7735 15988 7744
rect 15936 7701 15945 7735
rect 15945 7701 15979 7735
rect 15979 7701 15988 7735
rect 15936 7692 15988 7701
rect 3519 7590 3571 7642
rect 3583 7590 3635 7642
rect 3647 7590 3699 7642
rect 3711 7590 3763 7642
rect 3775 7590 3827 7642
rect 7337 7590 7389 7642
rect 7401 7590 7453 7642
rect 7465 7590 7517 7642
rect 7529 7590 7581 7642
rect 7593 7590 7645 7642
rect 11155 7590 11207 7642
rect 11219 7590 11271 7642
rect 11283 7590 11335 7642
rect 11347 7590 11399 7642
rect 11411 7590 11463 7642
rect 14973 7590 15025 7642
rect 15037 7590 15089 7642
rect 15101 7590 15153 7642
rect 15165 7590 15217 7642
rect 15229 7590 15281 7642
rect 2044 7488 2096 7540
rect 2136 7488 2188 7540
rect 2412 7531 2464 7540
rect 2412 7497 2421 7531
rect 2421 7497 2455 7531
rect 2455 7497 2464 7531
rect 2412 7488 2464 7497
rect 940 7420 992 7472
rect 1860 7420 1912 7472
rect 1952 7463 2004 7472
rect 1952 7429 1961 7463
rect 1961 7429 1995 7463
rect 1995 7429 2004 7463
rect 1952 7420 2004 7429
rect 3884 7488 3936 7540
rect 3976 7488 4028 7540
rect 4160 7488 4212 7540
rect 4896 7488 4948 7540
rect 5540 7488 5592 7540
rect 2872 7463 2924 7472
rect 2872 7429 2881 7463
rect 2881 7429 2915 7463
rect 2915 7429 2924 7463
rect 2872 7420 2924 7429
rect 1768 7395 1820 7404
rect 1768 7361 1777 7395
rect 1777 7361 1811 7395
rect 1811 7361 1820 7395
rect 1768 7352 1820 7361
rect 2504 7352 2556 7404
rect 2320 7284 2372 7336
rect 3332 7216 3384 7268
rect 3792 7352 3844 7404
rect 5908 7488 5960 7540
rect 6460 7488 6512 7540
rect 7564 7488 7616 7540
rect 4528 7352 4580 7404
rect 3976 7327 4028 7336
rect 3976 7293 3985 7327
rect 3985 7293 4019 7327
rect 4019 7293 4028 7327
rect 3976 7284 4028 7293
rect 4252 7284 4304 7336
rect 5448 7352 5500 7404
rect 5816 7352 5868 7404
rect 8760 7488 8812 7540
rect 9036 7488 9088 7540
rect 10048 7488 10100 7540
rect 8024 7420 8076 7472
rect 8300 7420 8352 7472
rect 8484 7420 8536 7472
rect 9496 7463 9548 7472
rect 7288 7395 7340 7404
rect 7288 7361 7297 7395
rect 7297 7361 7331 7395
rect 7331 7361 7340 7395
rect 7288 7352 7340 7361
rect 7564 7395 7616 7404
rect 7564 7361 7573 7395
rect 7573 7361 7607 7395
rect 7607 7361 7616 7395
rect 7564 7352 7616 7361
rect 9496 7429 9505 7463
rect 9505 7429 9539 7463
rect 9539 7429 9548 7463
rect 9496 7420 9548 7429
rect 12440 7531 12492 7540
rect 12440 7497 12465 7531
rect 12465 7497 12492 7531
rect 12440 7488 12492 7497
rect 12900 7488 12952 7540
rect 13176 7488 13228 7540
rect 13636 7531 13688 7540
rect 13636 7497 13645 7531
rect 13645 7497 13679 7531
rect 13679 7497 13688 7531
rect 13636 7488 13688 7497
rect 14372 7488 14424 7540
rect 14832 7488 14884 7540
rect 9312 7352 9364 7404
rect 10140 7395 10192 7404
rect 10140 7361 10149 7395
rect 10149 7361 10183 7395
rect 10183 7361 10192 7395
rect 10140 7352 10192 7361
rect 10876 7420 10928 7472
rect 12164 7420 12216 7472
rect 7012 7216 7064 7268
rect 7840 7216 7892 7268
rect 2780 7148 2832 7200
rect 3792 7148 3844 7200
rect 4068 7148 4120 7200
rect 4712 7148 4764 7200
rect 4804 7191 4856 7200
rect 4804 7157 4813 7191
rect 4813 7157 4847 7191
rect 4847 7157 4856 7191
rect 4804 7148 4856 7157
rect 4896 7148 4948 7200
rect 5632 7148 5684 7200
rect 5816 7148 5868 7200
rect 6184 7148 6236 7200
rect 6552 7191 6604 7200
rect 6552 7157 6561 7191
rect 6561 7157 6595 7191
rect 6595 7157 6604 7191
rect 6552 7148 6604 7157
rect 7288 7148 7340 7200
rect 8668 7148 8720 7200
rect 9680 7191 9732 7200
rect 9680 7157 9689 7191
rect 9689 7157 9723 7191
rect 9723 7157 9732 7191
rect 9680 7148 9732 7157
rect 10416 7148 10468 7200
rect 12808 7216 12860 7268
rect 13360 7216 13412 7268
rect 14464 7463 14516 7472
rect 14464 7429 14473 7463
rect 14473 7429 14507 7463
rect 14507 7429 14516 7463
rect 14464 7420 14516 7429
rect 12072 7148 12124 7200
rect 2859 7046 2911 7098
rect 2923 7046 2975 7098
rect 2987 7046 3039 7098
rect 3051 7046 3103 7098
rect 3115 7046 3167 7098
rect 6677 7046 6729 7098
rect 6741 7046 6793 7098
rect 6805 7046 6857 7098
rect 6869 7046 6921 7098
rect 6933 7046 6985 7098
rect 10495 7046 10547 7098
rect 10559 7046 10611 7098
rect 10623 7046 10675 7098
rect 10687 7046 10739 7098
rect 10751 7046 10803 7098
rect 14313 7046 14365 7098
rect 14377 7046 14429 7098
rect 14441 7046 14493 7098
rect 14505 7046 14557 7098
rect 14569 7046 14621 7098
rect 1860 6944 1912 6996
rect 3332 6944 3384 6996
rect 3976 6944 4028 6996
rect 5816 6944 5868 6996
rect 6092 6987 6144 6996
rect 6092 6953 6101 6987
rect 6101 6953 6135 6987
rect 6135 6953 6144 6987
rect 6092 6944 6144 6953
rect 6184 6944 6236 6996
rect 7748 6944 7800 6996
rect 10140 6944 10192 6996
rect 12072 6944 12124 6996
rect 2688 6876 2740 6928
rect 1768 6851 1820 6860
rect 1768 6817 1777 6851
rect 1777 6817 1811 6851
rect 1811 6817 1820 6851
rect 1768 6808 1820 6817
rect 2044 6808 2096 6860
rect 1860 6740 1912 6792
rect 1768 6672 1820 6724
rect 3884 6740 3936 6792
rect 3976 6740 4028 6792
rect 4160 6783 4212 6792
rect 4160 6749 4169 6783
rect 4169 6749 4203 6783
rect 4203 6749 4212 6783
rect 4160 6740 4212 6749
rect 4436 6740 4488 6792
rect 5540 6876 5592 6928
rect 6460 6876 6512 6928
rect 7564 6876 7616 6928
rect 8116 6876 8168 6928
rect 4712 6808 4764 6860
rect 4804 6740 4856 6792
rect 5356 6740 5408 6792
rect 5540 6783 5592 6792
rect 5540 6749 5549 6783
rect 5549 6749 5583 6783
rect 5583 6749 5592 6783
rect 5540 6740 5592 6749
rect 6368 6808 6420 6860
rect 6920 6851 6972 6860
rect 6920 6817 6943 6851
rect 6943 6817 6972 6851
rect 6920 6808 6972 6817
rect 5632 6715 5684 6724
rect 5632 6681 5641 6715
rect 5641 6681 5675 6715
rect 5675 6681 5684 6715
rect 5632 6672 5684 6681
rect 2688 6604 2740 6656
rect 3240 6604 3292 6656
rect 4528 6604 4580 6656
rect 5080 6647 5132 6656
rect 5080 6613 5089 6647
rect 5089 6613 5123 6647
rect 5123 6613 5132 6647
rect 5080 6604 5132 6613
rect 5264 6647 5316 6656
rect 5264 6613 5273 6647
rect 5273 6613 5307 6647
rect 5307 6613 5316 6647
rect 6828 6715 6880 6724
rect 6828 6681 6837 6715
rect 6837 6681 6871 6715
rect 6871 6681 6880 6715
rect 6828 6672 6880 6681
rect 8116 6783 8168 6792
rect 8116 6749 8125 6783
rect 8125 6749 8159 6783
rect 8159 6749 8168 6783
rect 8116 6740 8168 6749
rect 8576 6740 8628 6792
rect 9496 6783 9548 6792
rect 9496 6749 9505 6783
rect 9505 6749 9539 6783
rect 9539 6749 9548 6783
rect 9496 6740 9548 6749
rect 9680 6876 9732 6928
rect 10416 6740 10468 6792
rect 10876 6783 10928 6792
rect 10876 6749 10885 6783
rect 10885 6749 10919 6783
rect 10919 6749 10928 6783
rect 10876 6740 10928 6749
rect 8760 6672 8812 6724
rect 9312 6715 9364 6724
rect 9312 6681 9321 6715
rect 9321 6681 9355 6715
rect 9355 6681 9364 6715
rect 9312 6672 9364 6681
rect 5264 6604 5316 6613
rect 7012 6647 7064 6656
rect 7012 6613 7021 6647
rect 7021 6613 7055 6647
rect 7055 6613 7064 6647
rect 7012 6604 7064 6613
rect 8024 6604 8076 6656
rect 8300 6647 8352 6656
rect 8300 6613 8309 6647
rect 8309 6613 8343 6647
rect 8343 6613 8352 6647
rect 8300 6604 8352 6613
rect 11612 6604 11664 6656
rect 12256 6783 12308 6792
rect 12256 6749 12265 6783
rect 12265 6749 12299 6783
rect 12299 6749 12308 6783
rect 12256 6740 12308 6749
rect 3519 6502 3571 6554
rect 3583 6502 3635 6554
rect 3647 6502 3699 6554
rect 3711 6502 3763 6554
rect 3775 6502 3827 6554
rect 7337 6502 7389 6554
rect 7401 6502 7453 6554
rect 7465 6502 7517 6554
rect 7529 6502 7581 6554
rect 7593 6502 7645 6554
rect 11155 6502 11207 6554
rect 11219 6502 11271 6554
rect 11283 6502 11335 6554
rect 11347 6502 11399 6554
rect 11411 6502 11463 6554
rect 14973 6502 15025 6554
rect 15037 6502 15089 6554
rect 15101 6502 15153 6554
rect 15165 6502 15217 6554
rect 15229 6502 15281 6554
rect 2320 6400 2372 6452
rect 940 6264 992 6316
rect 1860 6264 1912 6316
rect 2320 6307 2372 6316
rect 2320 6273 2329 6307
rect 2329 6273 2363 6307
rect 2363 6273 2372 6307
rect 2320 6264 2372 6273
rect 4160 6400 4212 6452
rect 3884 6332 3936 6384
rect 4712 6400 4764 6452
rect 7012 6400 7064 6452
rect 7104 6400 7156 6452
rect 7932 6400 7984 6452
rect 8300 6400 8352 6452
rect 9036 6443 9088 6452
rect 9036 6409 9045 6443
rect 9045 6409 9079 6443
rect 9079 6409 9088 6443
rect 9036 6400 9088 6409
rect 12808 6443 12860 6452
rect 12808 6409 12817 6443
rect 12817 6409 12851 6443
rect 12851 6409 12860 6443
rect 12808 6400 12860 6409
rect 14740 6400 14792 6452
rect 4988 6375 5040 6384
rect 4988 6341 5029 6375
rect 5029 6341 5040 6375
rect 4988 6332 5040 6341
rect 6828 6332 6880 6384
rect 8852 6375 8904 6384
rect 8852 6341 8861 6375
rect 8861 6341 8895 6375
rect 8895 6341 8904 6375
rect 8852 6332 8904 6341
rect 1676 6239 1728 6248
rect 1676 6205 1685 6239
rect 1685 6205 1719 6239
rect 1719 6205 1728 6239
rect 1676 6196 1728 6205
rect 1952 6196 2004 6248
rect 3240 6196 3292 6248
rect 3976 6264 4028 6316
rect 4160 6196 4212 6248
rect 4528 6264 4580 6316
rect 5264 6196 5316 6248
rect 5356 6196 5408 6248
rect 5908 6307 5960 6316
rect 5908 6273 5917 6307
rect 5917 6273 5951 6307
rect 5951 6273 5960 6307
rect 5908 6264 5960 6273
rect 6184 6264 6236 6316
rect 6368 6307 6420 6316
rect 6368 6273 6377 6307
rect 6377 6273 6411 6307
rect 6411 6273 6420 6307
rect 6368 6264 6420 6273
rect 6460 6264 6512 6316
rect 6644 6307 6696 6316
rect 6644 6273 6653 6307
rect 6653 6273 6687 6307
rect 6687 6273 6696 6307
rect 6644 6264 6696 6273
rect 6736 6307 6788 6316
rect 6736 6273 6745 6307
rect 6745 6273 6779 6307
rect 6779 6273 6788 6307
rect 6736 6264 6788 6273
rect 7840 6307 7892 6316
rect 7840 6273 7849 6307
rect 7849 6273 7883 6307
rect 7883 6273 7892 6307
rect 7840 6264 7892 6273
rect 8024 6307 8076 6316
rect 8024 6273 8033 6307
rect 8033 6273 8067 6307
rect 8067 6273 8076 6307
rect 8024 6264 8076 6273
rect 10048 6332 10100 6384
rect 7472 6196 7524 6248
rect 9404 6264 9456 6316
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 12256 6264 12308 6316
rect 12900 6264 12952 6316
rect 13912 6307 13964 6316
rect 13912 6273 13921 6307
rect 13921 6273 13955 6307
rect 13955 6273 13964 6307
rect 13912 6264 13964 6273
rect 8668 6196 8720 6248
rect 9588 6196 9640 6248
rect 11612 6239 11664 6248
rect 11612 6205 11621 6239
rect 11621 6205 11655 6239
rect 11655 6205 11664 6239
rect 11612 6196 11664 6205
rect 12440 6239 12492 6248
rect 12440 6205 12449 6239
rect 12449 6205 12483 6239
rect 12483 6205 12492 6239
rect 12440 6196 12492 6205
rect 12992 6239 13044 6248
rect 12992 6205 13001 6239
rect 13001 6205 13035 6239
rect 13035 6205 13044 6239
rect 12992 6196 13044 6205
rect 2412 6060 2464 6112
rect 3424 6060 3476 6112
rect 3884 6060 3936 6112
rect 4436 6060 4488 6112
rect 6000 6128 6052 6180
rect 6644 6128 6696 6180
rect 11796 6128 11848 6180
rect 14556 6264 14608 6316
rect 14740 6264 14792 6316
rect 5816 6060 5868 6112
rect 7656 6103 7708 6112
rect 7656 6069 7665 6103
rect 7665 6069 7699 6103
rect 7699 6069 7708 6103
rect 7656 6060 7708 6069
rect 8484 6103 8536 6112
rect 8484 6069 8493 6103
rect 8493 6069 8527 6103
rect 8527 6069 8536 6103
rect 8484 6060 8536 6069
rect 9404 6060 9456 6112
rect 10048 6060 10100 6112
rect 11612 6060 11664 6112
rect 11980 6103 12032 6112
rect 11980 6069 11989 6103
rect 11989 6069 12023 6103
rect 12023 6069 12032 6103
rect 11980 6060 12032 6069
rect 14096 6060 14148 6112
rect 2859 5958 2911 6010
rect 2923 5958 2975 6010
rect 2987 5958 3039 6010
rect 3051 5958 3103 6010
rect 3115 5958 3167 6010
rect 6677 5958 6729 6010
rect 6741 5958 6793 6010
rect 6805 5958 6857 6010
rect 6869 5958 6921 6010
rect 6933 5958 6985 6010
rect 10495 5958 10547 6010
rect 10559 5958 10611 6010
rect 10623 5958 10675 6010
rect 10687 5958 10739 6010
rect 10751 5958 10803 6010
rect 14313 5958 14365 6010
rect 14377 5958 14429 6010
rect 14441 5958 14493 6010
rect 14505 5958 14557 6010
rect 14569 5958 14621 6010
rect 1676 5856 1728 5908
rect 3332 5856 3384 5908
rect 4988 5856 5040 5908
rect 6092 5856 6144 5908
rect 6552 5856 6604 5908
rect 7472 5856 7524 5908
rect 7932 5856 7984 5908
rect 8300 5856 8352 5908
rect 8576 5856 8628 5908
rect 9036 5856 9088 5908
rect 9404 5856 9456 5908
rect 11704 5856 11756 5908
rect 11980 5856 12032 5908
rect 5632 5788 5684 5840
rect 2320 5720 2372 5772
rect 1952 5695 2004 5704
rect 1952 5661 1961 5695
rect 1961 5661 1995 5695
rect 1995 5661 2004 5695
rect 1952 5652 2004 5661
rect 2044 5652 2096 5704
rect 2596 5763 2648 5772
rect 2596 5729 2605 5763
rect 2605 5729 2639 5763
rect 2639 5729 2648 5763
rect 2596 5720 2648 5729
rect 2688 5720 2740 5772
rect 5816 5720 5868 5772
rect 6368 5720 6420 5772
rect 1676 5584 1728 5636
rect 1768 5627 1820 5636
rect 1768 5593 1777 5627
rect 1777 5593 1811 5627
rect 1811 5593 1820 5627
rect 1768 5584 1820 5593
rect 3148 5652 3200 5704
rect 4160 5652 4212 5704
rect 4528 5695 4580 5704
rect 4528 5661 4540 5695
rect 4540 5661 4574 5695
rect 4574 5661 4580 5695
rect 4528 5652 4580 5661
rect 1860 5516 1912 5568
rect 2136 5559 2188 5568
rect 2136 5525 2145 5559
rect 2145 5525 2179 5559
rect 2179 5525 2188 5559
rect 2136 5516 2188 5525
rect 4436 5584 4488 5636
rect 4804 5695 4856 5704
rect 4804 5661 4813 5695
rect 4813 5661 4847 5695
rect 4847 5661 4856 5695
rect 4804 5652 4856 5661
rect 6000 5695 6052 5704
rect 6000 5661 6009 5695
rect 6009 5661 6043 5695
rect 6043 5661 6052 5695
rect 6000 5652 6052 5661
rect 6092 5695 6144 5704
rect 6092 5661 6101 5695
rect 6101 5661 6135 5695
rect 6135 5661 6144 5695
rect 6092 5652 6144 5661
rect 6184 5695 6236 5704
rect 6184 5661 6193 5695
rect 6193 5661 6227 5695
rect 6227 5661 6236 5695
rect 6184 5652 6236 5661
rect 6000 5516 6052 5568
rect 8024 5788 8076 5840
rect 8392 5720 8444 5772
rect 7656 5652 7708 5704
rect 7932 5652 7984 5704
rect 8484 5652 8536 5704
rect 8208 5559 8260 5568
rect 8208 5525 8217 5559
rect 8217 5525 8251 5559
rect 8251 5525 8260 5559
rect 8208 5516 8260 5525
rect 8300 5516 8352 5568
rect 8576 5516 8628 5568
rect 9588 5695 9640 5704
rect 9588 5661 9597 5695
rect 9597 5661 9631 5695
rect 9631 5661 9640 5695
rect 9588 5652 9640 5661
rect 11520 5788 11572 5840
rect 11612 5831 11664 5840
rect 11612 5797 11621 5831
rect 11621 5797 11655 5831
rect 11655 5797 11664 5831
rect 11612 5788 11664 5797
rect 12992 5856 13044 5908
rect 14648 5899 14700 5908
rect 14648 5865 14657 5899
rect 14657 5865 14691 5899
rect 14691 5865 14700 5899
rect 14648 5856 14700 5865
rect 14096 5720 14148 5772
rect 11796 5652 11848 5704
rect 12900 5652 12952 5704
rect 13360 5695 13412 5704
rect 13360 5661 13369 5695
rect 13369 5661 13403 5695
rect 13403 5661 13412 5695
rect 13360 5652 13412 5661
rect 13912 5652 13964 5704
rect 14740 5652 14792 5704
rect 9680 5516 9732 5568
rect 11612 5516 11664 5568
rect 12440 5516 12492 5568
rect 13176 5516 13228 5568
rect 16028 5516 16080 5568
rect 3519 5414 3571 5466
rect 3583 5414 3635 5466
rect 3647 5414 3699 5466
rect 3711 5414 3763 5466
rect 3775 5414 3827 5466
rect 7337 5414 7389 5466
rect 7401 5414 7453 5466
rect 7465 5414 7517 5466
rect 7529 5414 7581 5466
rect 7593 5414 7645 5466
rect 11155 5414 11207 5466
rect 11219 5414 11271 5466
rect 11283 5414 11335 5466
rect 11347 5414 11399 5466
rect 11411 5414 11463 5466
rect 14973 5414 15025 5466
rect 15037 5414 15089 5466
rect 15101 5414 15153 5466
rect 15165 5414 15217 5466
rect 15229 5414 15281 5466
rect 4344 5312 4396 5364
rect 4528 5312 4580 5364
rect 8392 5312 8444 5364
rect 8484 5312 8536 5364
rect 2504 5244 2556 5296
rect 2780 5244 2832 5296
rect 3148 5244 3200 5296
rect 1676 5176 1728 5228
rect 2596 5108 2648 5160
rect 3516 5108 3568 5160
rect 4252 5219 4304 5228
rect 4252 5185 4261 5219
rect 4261 5185 4295 5219
rect 4295 5185 4304 5219
rect 7840 5287 7892 5296
rect 7840 5253 7849 5287
rect 7849 5253 7883 5287
rect 7883 5253 7892 5287
rect 7840 5244 7892 5253
rect 7932 5287 7984 5296
rect 7932 5253 7941 5287
rect 7941 5253 7975 5287
rect 7975 5253 7984 5287
rect 7932 5244 7984 5253
rect 4252 5176 4304 5185
rect 5080 5176 5132 5228
rect 6368 5219 6420 5228
rect 6368 5185 6377 5219
rect 6377 5185 6411 5219
rect 6411 5185 6420 5219
rect 6368 5176 6420 5185
rect 5356 5151 5408 5160
rect 5356 5117 5365 5151
rect 5365 5117 5399 5151
rect 5399 5117 5408 5151
rect 5356 5108 5408 5117
rect 8300 5176 8352 5228
rect 8668 5176 8720 5228
rect 9680 5312 9732 5364
rect 13360 5312 13412 5364
rect 8392 5108 8444 5160
rect 11520 5287 11572 5296
rect 11520 5253 11529 5287
rect 11529 5253 11563 5287
rect 11563 5253 11572 5287
rect 11520 5244 11572 5253
rect 11704 5287 11756 5296
rect 11704 5253 11713 5287
rect 11713 5253 11747 5287
rect 11747 5253 11756 5287
rect 11704 5244 11756 5253
rect 9404 5040 9456 5092
rect 12992 5176 13044 5228
rect 13176 5219 13228 5228
rect 13176 5185 13185 5219
rect 13185 5185 13219 5219
rect 13219 5185 13228 5219
rect 13176 5176 13228 5185
rect 3976 5015 4028 5024
rect 3976 4981 3985 5015
rect 3985 4981 4019 5015
rect 4019 4981 4028 5015
rect 3976 4972 4028 4981
rect 4160 4972 4212 5024
rect 6092 4972 6144 5024
rect 8760 5015 8812 5024
rect 8760 4981 8769 5015
rect 8769 4981 8803 5015
rect 8803 4981 8812 5015
rect 8760 4972 8812 4981
rect 8944 5015 8996 5024
rect 8944 4981 8953 5015
rect 8953 4981 8987 5015
rect 8987 4981 8996 5015
rect 8944 4972 8996 4981
rect 10048 5015 10100 5024
rect 10048 4981 10057 5015
rect 10057 4981 10091 5015
rect 10091 4981 10100 5015
rect 10048 4972 10100 4981
rect 10416 5015 10468 5024
rect 10416 4981 10425 5015
rect 10425 4981 10459 5015
rect 10459 4981 10468 5015
rect 10416 4972 10468 4981
rect 10876 4972 10928 5024
rect 11244 4972 11296 5024
rect 11888 5015 11940 5024
rect 11888 4981 11897 5015
rect 11897 4981 11931 5015
rect 11931 4981 11940 5015
rect 11888 4972 11940 4981
rect 2859 4870 2911 4922
rect 2923 4870 2975 4922
rect 2987 4870 3039 4922
rect 3051 4870 3103 4922
rect 3115 4870 3167 4922
rect 6677 4870 6729 4922
rect 6741 4870 6793 4922
rect 6805 4870 6857 4922
rect 6869 4870 6921 4922
rect 6933 4870 6985 4922
rect 10495 4870 10547 4922
rect 10559 4870 10611 4922
rect 10623 4870 10675 4922
rect 10687 4870 10739 4922
rect 10751 4870 10803 4922
rect 14313 4870 14365 4922
rect 14377 4870 14429 4922
rect 14441 4870 14493 4922
rect 14505 4870 14557 4922
rect 14569 4870 14621 4922
rect 1768 4675 1820 4684
rect 1768 4641 1777 4675
rect 1777 4641 1811 4675
rect 1811 4641 1820 4675
rect 1768 4632 1820 4641
rect 940 4564 992 4616
rect 2136 4564 2188 4616
rect 2780 4632 2832 4684
rect 2412 4564 2464 4616
rect 3516 4768 3568 4820
rect 3976 4768 4028 4820
rect 6092 4700 6144 4752
rect 2596 4496 2648 4548
rect 4160 4607 4212 4616
rect 4160 4573 4169 4607
rect 4169 4573 4203 4607
rect 4203 4573 4212 4607
rect 4160 4564 4212 4573
rect 7012 4768 7064 4820
rect 10416 4768 10468 4820
rect 10876 4768 10928 4820
rect 11612 4768 11664 4820
rect 6368 4700 6420 4752
rect 7656 4632 7708 4684
rect 7104 4564 7156 4616
rect 7564 4564 7616 4616
rect 11244 4743 11296 4752
rect 11244 4709 11253 4743
rect 11253 4709 11287 4743
rect 11287 4709 11296 4743
rect 11244 4700 11296 4709
rect 11060 4632 11112 4684
rect 3332 4471 3384 4480
rect 3332 4437 3341 4471
rect 3341 4437 3375 4471
rect 3375 4437 3384 4471
rect 3332 4428 3384 4437
rect 4344 4471 4396 4480
rect 4344 4437 4353 4471
rect 4353 4437 4387 4471
rect 4387 4437 4396 4471
rect 4344 4428 4396 4437
rect 7564 4428 7616 4480
rect 3519 4326 3571 4378
rect 3583 4326 3635 4378
rect 3647 4326 3699 4378
rect 3711 4326 3763 4378
rect 3775 4326 3827 4378
rect 7337 4326 7389 4378
rect 7401 4326 7453 4378
rect 7465 4326 7517 4378
rect 7529 4326 7581 4378
rect 7593 4326 7645 4378
rect 11155 4326 11207 4378
rect 11219 4326 11271 4378
rect 11283 4326 11335 4378
rect 11347 4326 11399 4378
rect 11411 4326 11463 4378
rect 14973 4326 15025 4378
rect 15037 4326 15089 4378
rect 15101 4326 15153 4378
rect 15165 4326 15217 4378
rect 15229 4326 15281 4378
rect 1860 4224 1912 4276
rect 3884 4224 3936 4276
rect 4896 4224 4948 4276
rect 1032 4156 1084 4208
rect 2780 4199 2832 4208
rect 2780 4165 2789 4199
rect 2789 4165 2823 4199
rect 2823 4165 2832 4199
rect 2780 4156 2832 4165
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 1676 4131 1728 4140
rect 1676 4097 1685 4131
rect 1685 4097 1719 4131
rect 1719 4097 1728 4131
rect 1676 4088 1728 4097
rect 3332 4156 3384 4208
rect 4068 4088 4120 4140
rect 4344 4088 4396 4140
rect 7012 4088 7064 4140
rect 8944 4088 8996 4140
rect 3240 3952 3292 4004
rect 4252 4063 4304 4072
rect 4252 4029 4261 4063
rect 4261 4029 4295 4063
rect 4295 4029 4304 4063
rect 4252 4020 4304 4029
rect 7656 4020 7708 4072
rect 11060 4088 11112 4140
rect 11888 4088 11940 4140
rect 8300 3952 8352 4004
rect 3332 3884 3384 3936
rect 3976 3884 4028 3936
rect 4436 3927 4488 3936
rect 4436 3893 4445 3927
rect 4445 3893 4479 3927
rect 4479 3893 4488 3927
rect 4436 3884 4488 3893
rect 7196 3884 7248 3936
rect 8116 3884 8168 3936
rect 8944 3884 8996 3936
rect 9128 3927 9180 3936
rect 9128 3893 9137 3927
rect 9137 3893 9171 3927
rect 9171 3893 9180 3927
rect 9128 3884 9180 3893
rect 9680 3927 9732 3936
rect 9680 3893 9689 3927
rect 9689 3893 9723 3927
rect 9723 3893 9732 3927
rect 9680 3884 9732 3893
rect 12900 4131 12952 4140
rect 12900 4097 12909 4131
rect 12909 4097 12943 4131
rect 12943 4097 12952 4131
rect 12900 4088 12952 4097
rect 13728 4131 13780 4140
rect 13728 4097 13737 4131
rect 13737 4097 13771 4131
rect 13771 4097 13780 4131
rect 13728 4088 13780 4097
rect 14004 4131 14056 4140
rect 14004 4097 14013 4131
rect 14013 4097 14047 4131
rect 14047 4097 14056 4131
rect 14004 4088 14056 4097
rect 14096 4131 14148 4140
rect 14096 4097 14105 4131
rect 14105 4097 14139 4131
rect 14139 4097 14148 4131
rect 14096 4088 14148 4097
rect 14740 4088 14792 4140
rect 12532 3952 12584 4004
rect 12624 3884 12676 3936
rect 13544 3884 13596 3936
rect 2859 3782 2911 3834
rect 2923 3782 2975 3834
rect 2987 3782 3039 3834
rect 3051 3782 3103 3834
rect 3115 3782 3167 3834
rect 6677 3782 6729 3834
rect 6741 3782 6793 3834
rect 6805 3782 6857 3834
rect 6869 3782 6921 3834
rect 6933 3782 6985 3834
rect 10495 3782 10547 3834
rect 10559 3782 10611 3834
rect 10623 3782 10675 3834
rect 10687 3782 10739 3834
rect 10751 3782 10803 3834
rect 14313 3782 14365 3834
rect 14377 3782 14429 3834
rect 14441 3782 14493 3834
rect 14505 3782 14557 3834
rect 14569 3782 14621 3834
rect 5356 3680 5408 3732
rect 6276 3680 6328 3732
rect 7012 3680 7064 3732
rect 7840 3680 7892 3732
rect 8300 3680 8352 3732
rect 9128 3680 9180 3732
rect 9680 3680 9732 3732
rect 13728 3680 13780 3732
rect 14004 3680 14056 3732
rect 3424 3544 3476 3596
rect 4436 3544 4488 3596
rect 940 3476 992 3528
rect 6092 3544 6144 3596
rect 4620 3408 4672 3460
rect 6276 3476 6328 3528
rect 6736 3655 6788 3664
rect 6736 3621 6745 3655
rect 6745 3621 6779 3655
rect 6779 3621 6788 3655
rect 6736 3612 6788 3621
rect 6920 3612 6972 3664
rect 6368 3408 6420 3460
rect 4160 3383 4212 3392
rect 4160 3349 4169 3383
rect 4169 3349 4203 3383
rect 4203 3349 4212 3383
rect 4160 3340 4212 3349
rect 5632 3383 5684 3392
rect 5632 3349 5641 3383
rect 5641 3349 5675 3383
rect 5675 3349 5684 3383
rect 5632 3340 5684 3349
rect 5816 3340 5868 3392
rect 6552 3451 6604 3460
rect 6552 3417 6561 3451
rect 6561 3417 6595 3451
rect 6595 3417 6604 3451
rect 6552 3408 6604 3417
rect 8208 3476 8260 3528
rect 12624 3587 12676 3596
rect 12624 3553 12633 3587
rect 12633 3553 12667 3587
rect 12667 3553 12676 3587
rect 12624 3544 12676 3553
rect 12532 3476 12584 3528
rect 15936 3655 15988 3664
rect 15936 3621 15945 3655
rect 15945 3621 15979 3655
rect 15979 3621 15988 3655
rect 15936 3612 15988 3621
rect 13544 3519 13596 3528
rect 13544 3485 13553 3519
rect 13553 3485 13587 3519
rect 13587 3485 13596 3519
rect 13544 3476 13596 3485
rect 14096 3408 14148 3460
rect 7012 3340 7064 3392
rect 9312 3340 9364 3392
rect 13176 3340 13228 3392
rect 3519 3238 3571 3290
rect 3583 3238 3635 3290
rect 3647 3238 3699 3290
rect 3711 3238 3763 3290
rect 3775 3238 3827 3290
rect 7337 3238 7389 3290
rect 7401 3238 7453 3290
rect 7465 3238 7517 3290
rect 7529 3238 7581 3290
rect 7593 3238 7645 3290
rect 11155 3238 11207 3290
rect 11219 3238 11271 3290
rect 11283 3238 11335 3290
rect 11347 3238 11399 3290
rect 11411 3238 11463 3290
rect 14973 3238 15025 3290
rect 15037 3238 15089 3290
rect 15101 3238 15153 3290
rect 15165 3238 15217 3290
rect 15229 3238 15281 3290
rect 3332 3136 3384 3188
rect 4160 3136 4212 3188
rect 4620 3136 4672 3188
rect 5632 3136 5684 3188
rect 940 3000 992 3052
rect 1952 2975 2004 2984
rect 1952 2941 1961 2975
rect 1961 2941 1995 2975
rect 1995 2941 2004 2975
rect 1952 2932 2004 2941
rect 3976 2932 4028 2984
rect 5356 3000 5408 3052
rect 7012 3179 7064 3188
rect 7012 3145 7021 3179
rect 7021 3145 7055 3179
rect 7055 3145 7064 3179
rect 7012 3136 7064 3145
rect 7656 3111 7708 3120
rect 7656 3077 7665 3111
rect 7665 3077 7699 3111
rect 7699 3077 7708 3111
rect 7656 3068 7708 3077
rect 5816 3043 5868 3052
rect 5816 3009 5825 3043
rect 5825 3009 5859 3043
rect 5859 3009 5868 3043
rect 5816 3000 5868 3009
rect 6920 3043 6972 3052
rect 6920 3009 6929 3043
rect 6929 3009 6963 3043
rect 6963 3009 6972 3043
rect 6920 3000 6972 3009
rect 4344 2864 4396 2916
rect 7196 2932 7248 2984
rect 8208 3068 8260 3120
rect 8576 3136 8628 3188
rect 8484 3068 8536 3120
rect 7196 2839 7248 2848
rect 7196 2805 7205 2839
rect 7205 2805 7239 2839
rect 7239 2805 7248 2839
rect 7196 2796 7248 2805
rect 7748 2932 7800 2984
rect 8576 3043 8628 3052
rect 8576 3009 8585 3043
rect 8585 3009 8619 3043
rect 8619 3009 8628 3043
rect 8576 3000 8628 3009
rect 9312 3068 9364 3120
rect 8392 2864 8444 2916
rect 9772 3000 9824 3052
rect 9128 2932 9180 2984
rect 10416 2932 10468 2984
rect 11428 2932 11480 2984
rect 11612 2975 11664 2984
rect 11612 2941 11621 2975
rect 11621 2941 11655 2975
rect 11655 2941 11664 2975
rect 11612 2932 11664 2941
rect 12440 2864 12492 2916
rect 7932 2796 7984 2848
rect 8484 2839 8536 2848
rect 8484 2805 8493 2839
rect 8493 2805 8527 2839
rect 8527 2805 8536 2839
rect 8484 2796 8536 2805
rect 8576 2839 8628 2848
rect 8576 2805 8585 2839
rect 8585 2805 8619 2839
rect 8619 2805 8628 2839
rect 8576 2796 8628 2805
rect 10876 2839 10928 2848
rect 10876 2805 10885 2839
rect 10885 2805 10919 2839
rect 10919 2805 10928 2839
rect 10876 2796 10928 2805
rect 13176 2796 13228 2848
rect 2859 2694 2911 2746
rect 2923 2694 2975 2746
rect 2987 2694 3039 2746
rect 3051 2694 3103 2746
rect 3115 2694 3167 2746
rect 6677 2694 6729 2746
rect 6741 2694 6793 2746
rect 6805 2694 6857 2746
rect 6869 2694 6921 2746
rect 6933 2694 6985 2746
rect 10495 2694 10547 2746
rect 10559 2694 10611 2746
rect 10623 2694 10675 2746
rect 10687 2694 10739 2746
rect 10751 2694 10803 2746
rect 14313 2694 14365 2746
rect 14377 2694 14429 2746
rect 14441 2694 14493 2746
rect 14505 2694 14557 2746
rect 14569 2694 14621 2746
rect 7104 2592 7156 2644
rect 7748 2635 7800 2644
rect 7748 2601 7757 2635
rect 7757 2601 7791 2635
rect 7791 2601 7800 2635
rect 7748 2592 7800 2601
rect 8024 2635 8076 2644
rect 8024 2601 8033 2635
rect 8033 2601 8067 2635
rect 8067 2601 8076 2635
rect 8024 2592 8076 2601
rect 9404 2592 9456 2644
rect 10876 2592 10928 2644
rect 7196 2524 7248 2576
rect 4344 2388 4396 2440
rect 7196 2431 7248 2440
rect 7196 2397 7205 2431
rect 7205 2397 7239 2431
rect 7239 2397 7248 2431
rect 7196 2388 7248 2397
rect 8484 2456 8536 2508
rect 8576 2388 8628 2440
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 9956 2388 10008 2440
rect 10416 2388 10468 2440
rect 12440 2431 12492 2440
rect 12440 2397 12449 2431
rect 12449 2397 12483 2431
rect 12483 2397 12492 2431
rect 12440 2388 12492 2397
rect 4528 2252 4580 2304
rect 7748 2252 7800 2304
rect 8392 2295 8444 2304
rect 8392 2261 8401 2295
rect 8401 2261 8435 2295
rect 8435 2261 8444 2295
rect 8392 2252 8444 2261
rect 12348 2252 12400 2304
rect 3519 2150 3571 2202
rect 3583 2150 3635 2202
rect 3647 2150 3699 2202
rect 3711 2150 3763 2202
rect 3775 2150 3827 2202
rect 7337 2150 7389 2202
rect 7401 2150 7453 2202
rect 7465 2150 7517 2202
rect 7529 2150 7581 2202
rect 7593 2150 7645 2202
rect 11155 2150 11207 2202
rect 11219 2150 11271 2202
rect 11283 2150 11335 2202
rect 11347 2150 11399 2202
rect 11411 2150 11463 2202
rect 14973 2150 15025 2202
rect 15037 2150 15089 2202
rect 15101 2150 15153 2202
rect 15165 2150 15217 2202
rect 15229 2150 15281 2202
<< metal2 >>
rect 12254 18843 12310 19643
rect 13542 18986 13598 19643
rect 13542 18958 13768 18986
rect 13542 18843 13598 18958
rect 12268 17898 12296 18843
rect 12268 17870 12480 17898
rect 3519 17436 3827 17445
rect 3519 17434 3525 17436
rect 3581 17434 3605 17436
rect 3661 17434 3685 17436
rect 3741 17434 3765 17436
rect 3821 17434 3827 17436
rect 3581 17382 3583 17434
rect 3763 17382 3765 17434
rect 3519 17380 3525 17382
rect 3581 17380 3605 17382
rect 3661 17380 3685 17382
rect 3741 17380 3765 17382
rect 3821 17380 3827 17382
rect 3519 17371 3827 17380
rect 7337 17436 7645 17445
rect 7337 17434 7343 17436
rect 7399 17434 7423 17436
rect 7479 17434 7503 17436
rect 7559 17434 7583 17436
rect 7639 17434 7645 17436
rect 7399 17382 7401 17434
rect 7581 17382 7583 17434
rect 7337 17380 7343 17382
rect 7399 17380 7423 17382
rect 7479 17380 7503 17382
rect 7559 17380 7583 17382
rect 7639 17380 7645 17382
rect 7337 17371 7645 17380
rect 11155 17436 11463 17445
rect 11155 17434 11161 17436
rect 11217 17434 11241 17436
rect 11297 17434 11321 17436
rect 11377 17434 11401 17436
rect 11457 17434 11463 17436
rect 11217 17382 11219 17434
rect 11399 17382 11401 17434
rect 11155 17380 11161 17382
rect 11217 17380 11241 17382
rect 11297 17380 11321 17382
rect 11377 17380 11401 17382
rect 11457 17380 11463 17382
rect 11155 17371 11463 17380
rect 12452 17270 12480 17870
rect 13740 17354 13768 18958
rect 14830 18843 14886 19643
rect 13740 17338 13860 17354
rect 14844 17338 14872 18843
rect 14973 17436 15281 17445
rect 14973 17434 14979 17436
rect 15035 17434 15059 17436
rect 15115 17434 15139 17436
rect 15195 17434 15219 17436
rect 15275 17434 15281 17436
rect 15035 17382 15037 17434
rect 15217 17382 15219 17434
rect 14973 17380 14979 17382
rect 15035 17380 15059 17382
rect 15115 17380 15139 17382
rect 15195 17380 15219 17382
rect 15275 17380 15281 17382
rect 14973 17371 15281 17380
rect 13740 17332 13872 17338
rect 13740 17326 13820 17332
rect 13820 17274 13872 17280
rect 14832 17332 14884 17338
rect 14832 17274 14884 17280
rect 12440 17264 12492 17270
rect 12440 17206 12492 17212
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 7288 17196 7340 17202
rect 7288 17138 7340 17144
rect 8024 17196 8076 17202
rect 8024 17138 8076 17144
rect 10324 17196 10376 17202
rect 10324 17138 10376 17144
rect 10416 17196 10468 17202
rect 10416 17138 10468 17144
rect 12164 17196 12216 17202
rect 12164 17138 12216 17144
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 14188 17196 14240 17202
rect 14188 17138 14240 17144
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 2859 16892 3167 16901
rect 2859 16890 2865 16892
rect 2921 16890 2945 16892
rect 3001 16890 3025 16892
rect 3081 16890 3105 16892
rect 3161 16890 3167 16892
rect 2921 16838 2923 16890
rect 3103 16838 3105 16890
rect 2859 16836 2865 16838
rect 2921 16836 2945 16838
rect 3001 16836 3025 16838
rect 3081 16836 3105 16838
rect 3161 16836 3167 16838
rect 2859 16827 3167 16836
rect 6677 16892 6985 16901
rect 6677 16890 6683 16892
rect 6739 16890 6763 16892
rect 6819 16890 6843 16892
rect 6899 16890 6923 16892
rect 6979 16890 6985 16892
rect 6739 16838 6741 16890
rect 6921 16838 6923 16890
rect 6677 16836 6683 16838
rect 6739 16836 6763 16838
rect 6819 16836 6843 16838
rect 6899 16836 6923 16838
rect 6979 16836 6985 16838
rect 6677 16827 6985 16836
rect 7208 16794 7236 17138
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 6000 16584 6052 16590
rect 6000 16526 6052 16532
rect 7196 16584 7248 16590
rect 7300 16572 7328 17138
rect 7472 17060 7524 17066
rect 7472 17002 7524 17008
rect 7484 16794 7512 17002
rect 8036 16794 8064 17138
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 9048 16794 9076 16934
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 9036 16788 9088 16794
rect 9036 16730 9088 16736
rect 8036 16590 8064 16730
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 7248 16544 7328 16572
rect 7932 16584 7984 16590
rect 7196 16526 7248 16532
rect 7932 16526 7984 16532
rect 8024 16584 8076 16590
rect 8024 16526 8076 16532
rect 3519 16348 3827 16357
rect 3519 16346 3525 16348
rect 3581 16346 3605 16348
rect 3661 16346 3685 16348
rect 3741 16346 3765 16348
rect 3821 16346 3827 16348
rect 3581 16294 3583 16346
rect 3763 16294 3765 16346
rect 3519 16292 3525 16294
rect 3581 16292 3605 16294
rect 3661 16292 3685 16294
rect 3741 16292 3765 16294
rect 3821 16292 3827 16294
rect 3519 16283 3827 16292
rect 4160 16108 4212 16114
rect 4160 16050 4212 16056
rect 5632 16108 5684 16114
rect 5632 16050 5684 16056
rect 2859 15804 3167 15813
rect 2859 15802 2865 15804
rect 2921 15802 2945 15804
rect 3001 15802 3025 15804
rect 3081 15802 3105 15804
rect 3161 15802 3167 15804
rect 2921 15750 2923 15802
rect 3103 15750 3105 15802
rect 2859 15748 2865 15750
rect 2921 15748 2945 15750
rect 3001 15748 3025 15750
rect 3081 15748 3105 15750
rect 3161 15748 3167 15750
rect 2859 15739 3167 15748
rect 3519 15260 3827 15269
rect 3519 15258 3525 15260
rect 3581 15258 3605 15260
rect 3661 15258 3685 15260
rect 3741 15258 3765 15260
rect 3821 15258 3827 15260
rect 3581 15206 3583 15258
rect 3763 15206 3765 15258
rect 3519 15204 3525 15206
rect 3581 15204 3605 15206
rect 3661 15204 3685 15206
rect 3741 15204 3765 15206
rect 3821 15204 3827 15206
rect 3519 15195 3827 15204
rect 4172 15178 4200 16050
rect 3896 15150 4200 15178
rect 3896 15094 3924 15150
rect 3884 15088 3936 15094
rect 3884 15030 3936 15036
rect 2688 15020 2740 15026
rect 2688 14962 2740 14968
rect 2136 14816 2188 14822
rect 2136 14758 2188 14764
rect 938 14376 994 14385
rect 938 14311 940 14320
rect 992 14311 994 14320
rect 940 14282 992 14288
rect 1400 14272 1452 14278
rect 1400 14214 1452 14220
rect 1412 14006 1440 14214
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 1400 14000 1452 14006
rect 1400 13942 1452 13948
rect 1964 13870 1992 14010
rect 1952 13864 2004 13870
rect 2004 13812 2084 13818
rect 1952 13806 2084 13812
rect 1964 13790 2084 13806
rect 1860 13728 1912 13734
rect 1860 13670 1912 13676
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1872 13394 1900 13670
rect 1860 13388 1912 13394
rect 1860 13330 1912 13336
rect 940 13320 992 13326
rect 940 13262 992 13268
rect 952 13025 980 13262
rect 1964 13258 1992 13670
rect 1952 13252 2004 13258
rect 1952 13194 2004 13200
rect 938 13016 994 13025
rect 938 12951 994 12960
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 12345 1440 12786
rect 1860 12776 1912 12782
rect 1860 12718 1912 12724
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1398 12336 1454 12345
rect 1398 12271 1454 12280
rect 1688 12238 1716 12582
rect 1676 12232 1728 12238
rect 1676 12174 1728 12180
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1412 10985 1440 11086
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 940 10668 992 10674
rect 940 10610 992 10616
rect 952 10305 980 10610
rect 938 10296 994 10305
rect 938 10231 994 10240
rect 1492 9920 1544 9926
rect 1492 9862 1544 9868
rect 1504 9625 1532 9862
rect 1490 9616 1546 9625
rect 1688 9586 1716 12174
rect 1490 9551 1546 9560
rect 1676 9580 1728 9586
rect 1676 9522 1728 9528
rect 938 8936 994 8945
rect 938 8871 940 8880
rect 992 8871 994 8880
rect 1768 8900 1820 8906
rect 940 8842 992 8848
rect 1768 8842 1820 8848
rect 1780 8090 1808 8842
rect 1768 8084 1820 8090
rect 1768 8026 1820 8032
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 938 7576 994 7585
rect 938 7511 994 7520
rect 952 7478 980 7511
rect 940 7472 992 7478
rect 940 7414 992 7420
rect 1780 7410 1808 7686
rect 1872 7478 1900 12718
rect 1964 12170 1992 13194
rect 2056 12782 2084 13790
rect 2148 13394 2176 14758
rect 2596 14340 2648 14346
rect 2596 14282 2648 14288
rect 2228 14272 2280 14278
rect 2228 14214 2280 14220
rect 2240 14074 2268 14214
rect 2228 14068 2280 14074
rect 2228 14010 2280 14016
rect 2240 13938 2268 14010
rect 2504 14000 2556 14006
rect 2608 13988 2636 14282
rect 2700 14278 2728 14962
rect 3792 14952 3844 14958
rect 3792 14894 3844 14900
rect 2859 14716 3167 14725
rect 2859 14714 2865 14716
rect 2921 14714 2945 14716
rect 3001 14714 3025 14716
rect 3081 14714 3105 14716
rect 3161 14714 3167 14716
rect 2921 14662 2923 14714
rect 3103 14662 3105 14714
rect 2859 14660 2865 14662
rect 2921 14660 2945 14662
rect 3001 14660 3025 14662
rect 3081 14660 3105 14662
rect 3161 14660 3167 14662
rect 2859 14651 3167 14660
rect 3332 14544 3384 14550
rect 3332 14486 3384 14492
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 2780 14340 2832 14346
rect 2780 14282 2832 14288
rect 2688 14272 2740 14278
rect 2688 14214 2740 14220
rect 2556 13960 2636 13988
rect 2504 13942 2556 13948
rect 2228 13932 2280 13938
rect 2280 13892 2360 13920
rect 2228 13874 2280 13880
rect 2136 13388 2188 13394
rect 2136 13330 2188 13336
rect 2228 13320 2280 13326
rect 2228 13262 2280 13268
rect 2044 12776 2096 12782
rect 2044 12718 2096 12724
rect 2240 12646 2268 13262
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 2044 12436 2096 12442
rect 2332 12434 2360 13892
rect 2608 13530 2636 13960
rect 2688 13864 2740 13870
rect 2688 13806 2740 13812
rect 2596 13524 2648 13530
rect 2596 13466 2648 13472
rect 2504 13252 2556 13258
rect 2504 13194 2556 13200
rect 2412 13184 2464 13190
rect 2412 13126 2464 13132
rect 2096 12406 2360 12434
rect 2044 12378 2096 12384
rect 1952 12164 2004 12170
rect 1952 12106 2004 12112
rect 2228 12164 2280 12170
rect 2228 12106 2280 12112
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 1964 8090 1992 8366
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 2056 8022 2084 8366
rect 2044 8016 2096 8022
rect 2044 7958 2096 7964
rect 2044 7812 2096 7818
rect 2044 7754 2096 7760
rect 2056 7546 2084 7754
rect 2148 7546 2176 8434
rect 2240 8022 2268 12106
rect 2424 10742 2452 13126
rect 2516 12986 2544 13194
rect 2700 12986 2728 13806
rect 2792 13802 2820 14282
rect 3252 14074 3280 14350
rect 3240 14068 3292 14074
rect 3240 14010 3292 14016
rect 3344 13920 3372 14486
rect 3804 14482 3832 14894
rect 3896 14482 3924 15030
rect 5644 15026 5672 16050
rect 6012 15978 6040 16526
rect 6552 16516 6604 16522
rect 6552 16458 6604 16464
rect 6460 16448 6512 16454
rect 6460 16390 6512 16396
rect 6472 15978 6500 16390
rect 6000 15972 6052 15978
rect 6000 15914 6052 15920
rect 6460 15972 6512 15978
rect 6460 15914 6512 15920
rect 6012 15706 6040 15914
rect 6000 15700 6052 15706
rect 6000 15642 6052 15648
rect 6472 15638 6500 15914
rect 6460 15632 6512 15638
rect 6460 15574 6512 15580
rect 6564 15314 6592 16458
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 7104 16108 7156 16114
rect 7104 16050 7156 16056
rect 6840 15994 6868 16050
rect 6840 15966 7052 15994
rect 6677 15804 6985 15813
rect 6677 15802 6683 15804
rect 6739 15802 6763 15804
rect 6819 15802 6843 15804
rect 6899 15802 6923 15804
rect 6979 15802 6985 15804
rect 6739 15750 6741 15802
rect 6921 15750 6923 15802
rect 6677 15748 6683 15750
rect 6739 15748 6763 15750
rect 6819 15748 6843 15750
rect 6899 15748 6923 15750
rect 6979 15748 6985 15750
rect 6677 15739 6985 15748
rect 7024 15502 7052 15966
rect 7116 15502 7144 16050
rect 7208 15706 7236 16526
rect 7748 16448 7800 16454
rect 7748 16390 7800 16396
rect 7337 16348 7645 16357
rect 7337 16346 7343 16348
rect 7399 16346 7423 16348
rect 7479 16346 7503 16348
rect 7559 16346 7583 16348
rect 7639 16346 7645 16348
rect 7399 16294 7401 16346
rect 7581 16294 7583 16346
rect 7337 16292 7343 16294
rect 7399 16292 7423 16294
rect 7479 16292 7503 16294
rect 7559 16292 7583 16294
rect 7639 16292 7645 16294
rect 7337 16283 7645 16292
rect 7760 16250 7788 16390
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 7472 16176 7524 16182
rect 7472 16118 7524 16124
rect 7484 15706 7512 16118
rect 7944 15910 7972 16526
rect 8220 16182 8248 16594
rect 8944 16584 8996 16590
rect 8944 16526 8996 16532
rect 8208 16176 8260 16182
rect 8208 16118 8260 16124
rect 7748 15904 7800 15910
rect 7748 15846 7800 15852
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7012 15496 7064 15502
rect 7012 15438 7064 15444
rect 7104 15496 7156 15502
rect 7104 15438 7156 15444
rect 6644 15360 6696 15366
rect 6564 15308 6644 15314
rect 6564 15302 6696 15308
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 6564 15286 6684 15302
rect 6564 15162 6592 15286
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 4252 15020 4304 15026
rect 4252 14962 4304 14968
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 5632 15020 5684 15026
rect 5632 14962 5684 14968
rect 4068 14612 4120 14618
rect 4172 14600 4200 14962
rect 4120 14572 4200 14600
rect 4068 14554 4120 14560
rect 3516 14476 3568 14482
rect 3516 14418 3568 14424
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 3884 14476 3936 14482
rect 3884 14418 3936 14424
rect 3424 14340 3476 14346
rect 3424 14282 3476 14288
rect 3436 14074 3464 14282
rect 3528 14260 3556 14418
rect 4172 14414 4200 14572
rect 4264 14482 4292 14962
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 3608 14272 3660 14278
rect 3528 14232 3608 14260
rect 3608 14214 3660 14220
rect 3519 14172 3827 14181
rect 3519 14170 3525 14172
rect 3581 14170 3605 14172
rect 3661 14170 3685 14172
rect 3741 14170 3765 14172
rect 3821 14170 3827 14172
rect 3581 14118 3583 14170
rect 3763 14118 3765 14170
rect 3519 14116 3525 14118
rect 3581 14116 3605 14118
rect 3661 14116 3685 14118
rect 3741 14116 3765 14118
rect 3821 14116 3827 14118
rect 3519 14107 3827 14116
rect 3988 14074 4016 14350
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 4264 13938 4292 14418
rect 5184 14414 5212 14758
rect 5276 14618 5304 14962
rect 6552 14952 6604 14958
rect 6552 14894 6604 14900
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 5908 14408 5960 14414
rect 5908 14350 5960 14356
rect 3424 13932 3476 13938
rect 3344 13892 3424 13920
rect 3424 13874 3476 13880
rect 4252 13932 4304 13938
rect 4252 13874 4304 13880
rect 2780 13796 2832 13802
rect 2780 13738 2832 13744
rect 2792 13530 2820 13738
rect 4160 13728 4212 13734
rect 4160 13670 4212 13676
rect 2859 13628 3167 13637
rect 2859 13626 2865 13628
rect 2921 13626 2945 13628
rect 3001 13626 3025 13628
rect 3081 13626 3105 13628
rect 3161 13626 3167 13628
rect 2921 13574 2923 13626
rect 3103 13574 3105 13626
rect 2859 13572 2865 13574
rect 2921 13572 2945 13574
rect 3001 13572 3025 13574
rect 3081 13572 3105 13574
rect 3161 13572 3167 13574
rect 2859 13563 3167 13572
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 4172 13326 4200 13670
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 3252 12986 3280 13262
rect 3519 13084 3827 13093
rect 3519 13082 3525 13084
rect 3581 13082 3605 13084
rect 3661 13082 3685 13084
rect 3741 13082 3765 13084
rect 3821 13082 3827 13084
rect 3581 13030 3583 13082
rect 3763 13030 3765 13082
rect 3519 13028 3525 13030
rect 3581 13028 3605 13030
rect 3661 13028 3685 13030
rect 3741 13028 3765 13030
rect 3821 13028 3827 13030
rect 3519 13019 3827 13028
rect 2504 12980 2556 12986
rect 2504 12922 2556 12928
rect 2688 12980 2740 12986
rect 2688 12922 2740 12928
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 2700 12434 2728 12922
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 2859 12540 3167 12549
rect 2859 12538 2865 12540
rect 2921 12538 2945 12540
rect 3001 12538 3025 12540
rect 3081 12538 3105 12540
rect 3161 12538 3167 12540
rect 2921 12486 2923 12538
rect 3103 12486 3105 12538
rect 2859 12484 2865 12486
rect 2921 12484 2945 12486
rect 3001 12484 3025 12486
rect 3081 12484 3105 12486
rect 3161 12484 3167 12486
rect 2859 12475 3167 12484
rect 2516 12406 2728 12434
rect 2516 12238 2544 12406
rect 4264 12238 4292 12582
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 4252 12232 4304 12238
rect 4252 12174 4304 12180
rect 3240 12164 3292 12170
rect 3240 12106 3292 12112
rect 3252 11898 3280 12106
rect 3436 11898 3464 12174
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 3519 11996 3827 12005
rect 3519 11994 3525 11996
rect 3581 11994 3605 11996
rect 3661 11994 3685 11996
rect 3741 11994 3765 11996
rect 3821 11994 3827 11996
rect 3581 11942 3583 11994
rect 3763 11942 3765 11994
rect 3519 11940 3525 11942
rect 3581 11940 3605 11942
rect 3661 11940 3685 11942
rect 3741 11940 3765 11942
rect 3821 11940 3827 11942
rect 3519 11931 3827 11940
rect 4080 11898 4108 12038
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3424 11892 3476 11898
rect 3424 11834 3476 11840
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 4172 11762 4200 12174
rect 4264 11830 4292 12174
rect 4252 11824 4304 11830
rect 4252 11766 4304 11772
rect 4160 11756 4212 11762
rect 4160 11698 4212 11704
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 2859 11452 3167 11461
rect 2859 11450 2865 11452
rect 2921 11450 2945 11452
rect 3001 11450 3025 11452
rect 3081 11450 3105 11452
rect 3161 11450 3167 11452
rect 2921 11398 2923 11450
rect 3103 11398 3105 11450
rect 2859 11396 2865 11398
rect 2921 11396 2945 11398
rect 3001 11396 3025 11398
rect 3081 11396 3105 11398
rect 3161 11396 3167 11398
rect 2859 11387 3167 11396
rect 3519 10908 3827 10917
rect 3519 10906 3525 10908
rect 3581 10906 3605 10908
rect 3661 10906 3685 10908
rect 3741 10906 3765 10908
rect 3821 10906 3827 10908
rect 3581 10854 3583 10906
rect 3763 10854 3765 10906
rect 3519 10852 3525 10854
rect 3581 10852 3605 10854
rect 3661 10852 3685 10854
rect 3741 10852 3765 10854
rect 3821 10852 3827 10854
rect 3519 10843 3827 10852
rect 3896 10810 3924 11494
rect 4172 10810 4200 11698
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 2412 10736 2464 10742
rect 2412 10678 2464 10684
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2424 10266 2452 10542
rect 4436 10532 4488 10538
rect 4436 10474 4488 10480
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3608 10464 3660 10470
rect 3608 10406 3660 10412
rect 3884 10464 3936 10470
rect 3884 10406 3936 10412
rect 4344 10464 4396 10470
rect 4344 10406 4396 10412
rect 2859 10364 3167 10373
rect 2859 10362 2865 10364
rect 2921 10362 2945 10364
rect 3001 10362 3025 10364
rect 3081 10362 3105 10364
rect 3161 10362 3167 10364
rect 2921 10310 2923 10362
rect 3103 10310 3105 10362
rect 2859 10308 2865 10310
rect 2921 10308 2945 10310
rect 3001 10308 3025 10310
rect 3081 10308 3105 10310
rect 3161 10308 3167 10310
rect 2859 10299 3167 10308
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 3252 9722 3280 9998
rect 3436 9722 3464 10406
rect 3620 10198 3648 10406
rect 3896 10266 3924 10406
rect 3884 10260 3936 10266
rect 3884 10202 3936 10208
rect 4356 10198 4384 10406
rect 3608 10192 3660 10198
rect 3608 10134 3660 10140
rect 4344 10192 4396 10198
rect 4344 10134 4396 10140
rect 4448 10062 4476 10474
rect 4436 10056 4488 10062
rect 4436 9998 4488 10004
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 3519 9820 3827 9829
rect 3519 9818 3525 9820
rect 3581 9818 3605 9820
rect 3661 9818 3685 9820
rect 3741 9818 3765 9820
rect 3821 9818 3827 9820
rect 3581 9766 3583 9818
rect 3763 9766 3765 9818
rect 3519 9764 3525 9766
rect 3581 9764 3605 9766
rect 3661 9764 3685 9766
rect 3741 9764 3765 9766
rect 3821 9764 3827 9766
rect 3519 9755 3827 9764
rect 3240 9716 3292 9722
rect 3240 9658 3292 9664
rect 3424 9716 3476 9722
rect 3424 9658 3476 9664
rect 3252 9602 3280 9658
rect 3252 9586 3372 9602
rect 3252 9580 3384 9586
rect 3252 9574 3332 9580
rect 3332 9522 3384 9528
rect 3884 9376 3936 9382
rect 3884 9318 3936 9324
rect 2859 9276 3167 9285
rect 2859 9274 2865 9276
rect 2921 9274 2945 9276
rect 3001 9274 3025 9276
rect 3081 9274 3105 9276
rect 3161 9274 3167 9276
rect 2921 9222 2923 9274
rect 3103 9222 3105 9274
rect 2859 9220 2865 9222
rect 2921 9220 2945 9222
rect 3001 9220 3025 9222
rect 3081 9220 3105 9222
rect 3161 9220 3167 9222
rect 2859 9211 3167 9220
rect 3519 8732 3827 8741
rect 3519 8730 3525 8732
rect 3581 8730 3605 8732
rect 3661 8730 3685 8732
rect 3741 8730 3765 8732
rect 3821 8730 3827 8732
rect 3581 8678 3583 8730
rect 3763 8678 3765 8730
rect 3519 8676 3525 8678
rect 3581 8676 3605 8678
rect 3661 8676 3685 8678
rect 3741 8676 3765 8678
rect 3821 8676 3827 8678
rect 3519 8667 3827 8676
rect 3896 8634 3924 9318
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 2412 8288 2464 8294
rect 2412 8230 2464 8236
rect 2228 8016 2280 8022
rect 2228 7958 2280 7964
rect 2240 7886 2268 7958
rect 2424 7954 2452 8230
rect 2608 8090 2636 8434
rect 2780 8356 2832 8362
rect 2780 8298 2832 8304
rect 2686 8256 2742 8265
rect 2792 8242 2820 8298
rect 2742 8214 2820 8242
rect 2686 8191 2742 8200
rect 2859 8188 3167 8197
rect 2859 8186 2865 8188
rect 2921 8186 2945 8188
rect 3001 8186 3025 8188
rect 3081 8186 3105 8188
rect 3161 8186 3167 8188
rect 2921 8134 2923 8186
rect 3103 8134 3105 8186
rect 2859 8132 2865 8134
rect 2921 8132 2945 8134
rect 3001 8132 3025 8134
rect 3081 8132 3105 8134
rect 3161 8132 3167 8134
rect 2859 8123 3167 8132
rect 2596 8084 2648 8090
rect 2648 8044 2820 8072
rect 2596 8026 2648 8032
rect 2412 7948 2464 7954
rect 2412 7890 2464 7896
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 1860 7472 1912 7478
rect 1860 7414 1912 7420
rect 1952 7472 2004 7478
rect 2240 7426 2268 7822
rect 2424 7546 2452 7890
rect 2596 7880 2648 7886
rect 2502 7848 2558 7857
rect 2648 7840 2728 7868
rect 2596 7822 2648 7828
rect 2502 7783 2558 7792
rect 2516 7732 2544 7783
rect 2596 7744 2648 7750
rect 2516 7704 2596 7732
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2004 7420 2268 7426
rect 1952 7414 2268 7420
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 938 6896 994 6905
rect 1780 6866 1808 7346
rect 1872 7002 1900 7414
rect 1964 7398 2268 7414
rect 2516 7410 2544 7704
rect 2596 7686 2648 7692
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2320 7336 2372 7342
rect 2320 7278 2372 7284
rect 1860 6996 1912 7002
rect 1860 6938 1912 6944
rect 938 6831 994 6840
rect 1768 6860 1820 6866
rect 952 6322 980 6831
rect 1768 6802 1820 6808
rect 2044 6860 2096 6866
rect 2044 6802 2096 6808
rect 1860 6792 1912 6798
rect 1860 6734 1912 6740
rect 1768 6724 1820 6730
rect 1768 6666 1820 6672
rect 940 6316 992 6322
rect 940 6258 992 6264
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1688 5914 1716 6190
rect 1676 5908 1728 5914
rect 1676 5850 1728 5856
rect 1780 5642 1808 6666
rect 1872 6322 1900 6734
rect 1860 6316 1912 6322
rect 1860 6258 1912 6264
rect 1676 5636 1728 5642
rect 1676 5578 1728 5584
rect 1768 5636 1820 5642
rect 1768 5578 1820 5584
rect 938 5536 994 5545
rect 938 5471 994 5480
rect 952 4622 980 5471
rect 1688 5234 1716 5578
rect 1676 5228 1728 5234
rect 1676 5170 1728 5176
rect 1398 4720 1454 4729
rect 1398 4655 1454 4664
rect 940 4616 992 4622
rect 940 4558 992 4564
rect 1032 4208 1084 4214
rect 1030 4176 1032 4185
rect 1084 4176 1086 4185
rect 1412 4146 1440 4655
rect 1688 4146 1716 5170
rect 1780 4690 1808 5578
rect 1872 5574 1900 6258
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 1964 5710 1992 6190
rect 2056 5710 2084 6802
rect 2332 6458 2360 7278
rect 2320 6452 2372 6458
rect 2320 6394 2372 6400
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2332 5778 2360 6258
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2320 5772 2372 5778
rect 2320 5714 2372 5720
rect 1952 5704 2004 5710
rect 1952 5646 2004 5652
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 1860 5568 1912 5574
rect 1860 5510 1912 5516
rect 1768 4684 1820 4690
rect 1768 4626 1820 4632
rect 1872 4282 1900 5510
rect 1860 4276 1912 4282
rect 1860 4218 1912 4224
rect 1030 4111 1086 4120
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 940 3528 992 3534
rect 938 3496 940 3505
rect 992 3496 994 3505
rect 938 3431 994 3440
rect 940 3052 992 3058
rect 940 2994 992 3000
rect 952 2825 980 2994
rect 1964 2990 1992 5646
rect 2136 5568 2188 5574
rect 2136 5510 2188 5516
rect 2148 4622 2176 5510
rect 2424 4622 2452 6054
rect 2516 5302 2544 7346
rect 2700 6934 2728 7840
rect 2792 7206 2820 8044
rect 3436 7954 3464 8434
rect 3424 7948 3476 7954
rect 3424 7890 3476 7896
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 2884 7478 2912 7686
rect 2872 7472 2924 7478
rect 2872 7414 2924 7420
rect 3344 7274 3372 7822
rect 3528 7732 3556 8570
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 3608 7948 3660 7954
rect 3608 7890 3660 7896
rect 3620 7750 3648 7890
rect 3436 7704 3556 7732
rect 3608 7744 3660 7750
rect 3332 7268 3384 7274
rect 3332 7210 3384 7216
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2859 7100 3167 7109
rect 2859 7098 2865 7100
rect 2921 7098 2945 7100
rect 3001 7098 3025 7100
rect 3081 7098 3105 7100
rect 3161 7098 3167 7100
rect 2921 7046 2923 7098
rect 3103 7046 3105 7098
rect 2859 7044 2865 7046
rect 2921 7044 2945 7046
rect 3001 7044 3025 7046
rect 3081 7044 3105 7046
rect 3161 7044 3167 7046
rect 2859 7035 3167 7044
rect 3332 6996 3384 7002
rect 3332 6938 3384 6944
rect 2688 6928 2740 6934
rect 2688 6870 2740 6876
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 2700 5778 2728 6598
rect 3252 6254 3280 6598
rect 3240 6248 3292 6254
rect 2778 6216 2834 6225
rect 3240 6190 3292 6196
rect 2778 6151 2834 6160
rect 2596 5772 2648 5778
rect 2596 5714 2648 5720
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2504 5296 2556 5302
rect 2504 5238 2556 5244
rect 2608 5166 2636 5714
rect 2792 5302 2820 6151
rect 2859 6012 3167 6021
rect 2859 6010 2865 6012
rect 2921 6010 2945 6012
rect 3001 6010 3025 6012
rect 3081 6010 3105 6012
rect 3161 6010 3167 6012
rect 2921 5958 2923 6010
rect 3103 5958 3105 6010
rect 2859 5956 2865 5958
rect 2921 5956 2945 5958
rect 3001 5956 3025 5958
rect 3081 5956 3105 5958
rect 3161 5956 3167 5958
rect 2859 5947 3167 5956
rect 3252 5794 3280 6190
rect 3344 5914 3372 6938
rect 3436 6202 3464 7704
rect 3608 7686 3660 7692
rect 3519 7644 3827 7653
rect 3519 7642 3525 7644
rect 3581 7642 3605 7644
rect 3661 7642 3685 7644
rect 3741 7642 3765 7644
rect 3821 7642 3827 7644
rect 3581 7590 3583 7642
rect 3763 7590 3765 7642
rect 3519 7588 3525 7590
rect 3581 7588 3605 7590
rect 3661 7588 3685 7590
rect 3741 7588 3765 7590
rect 3821 7588 3827 7590
rect 3519 7579 3827 7588
rect 3896 7546 3924 8434
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3988 7546 4016 7686
rect 3884 7540 3936 7546
rect 3884 7482 3936 7488
rect 3976 7540 4028 7546
rect 3976 7482 4028 7488
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 3804 7206 3832 7346
rect 3792 7200 3844 7206
rect 3792 7142 3844 7148
rect 3896 6798 3924 7482
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 3988 7002 4016 7278
rect 4080 7206 4108 8434
rect 4172 7546 4200 9862
rect 4540 9654 4568 14350
rect 4988 14272 5040 14278
rect 4988 14214 5040 14220
rect 5080 14272 5132 14278
rect 5080 14214 5132 14220
rect 5000 13870 5028 14214
rect 5092 13938 5120 14214
rect 5184 14074 5212 14350
rect 5920 14074 5948 14350
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 4988 13864 5040 13870
rect 4988 13806 5040 13812
rect 4896 13184 4948 13190
rect 4896 13126 4948 13132
rect 4908 12986 4936 13126
rect 5000 12986 5028 13806
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 5092 12442 5120 13874
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 5264 13796 5316 13802
rect 5264 13738 5316 13744
rect 5276 13530 5304 13738
rect 5368 13530 5396 13806
rect 6564 13802 6592 14894
rect 7024 14822 7052 15302
rect 7116 15026 7144 15438
rect 7196 15428 7248 15434
rect 7196 15370 7248 15376
rect 7208 15094 7236 15370
rect 7337 15260 7645 15269
rect 7337 15258 7343 15260
rect 7399 15258 7423 15260
rect 7479 15258 7503 15260
rect 7559 15258 7583 15260
rect 7639 15258 7645 15260
rect 7399 15206 7401 15258
rect 7581 15206 7583 15258
rect 7337 15204 7343 15206
rect 7399 15204 7423 15206
rect 7479 15204 7503 15206
rect 7559 15204 7583 15206
rect 7639 15204 7645 15206
rect 7337 15195 7645 15204
rect 7196 15088 7248 15094
rect 7196 15030 7248 15036
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 7196 14816 7248 14822
rect 7196 14758 7248 14764
rect 6677 14716 6985 14725
rect 6677 14714 6683 14716
rect 6739 14714 6763 14716
rect 6819 14714 6843 14716
rect 6899 14714 6923 14716
rect 6979 14714 6985 14716
rect 6739 14662 6741 14714
rect 6921 14662 6923 14714
rect 6677 14660 6683 14662
rect 6739 14660 6763 14662
rect 6819 14660 6843 14662
rect 6899 14660 6923 14662
rect 6979 14660 6985 14662
rect 6677 14651 6985 14660
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6748 14074 6776 14214
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6552 13796 6604 13802
rect 6552 13738 6604 13744
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5908 13320 5960 13326
rect 5908 13262 5960 13268
rect 5552 12986 5580 13262
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5736 12442 5764 12786
rect 5920 12442 5948 13262
rect 5080 12436 5132 12442
rect 5080 12378 5132 12384
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4724 11898 4752 12174
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 5736 10810 5764 12378
rect 6012 12238 6040 13670
rect 6677 13628 6985 13637
rect 6677 13626 6683 13628
rect 6739 13626 6763 13628
rect 6819 13626 6843 13628
rect 6899 13626 6923 13628
rect 6979 13626 6985 13628
rect 6739 13574 6741 13626
rect 6921 13574 6923 13626
rect 6677 13572 6683 13574
rect 6739 13572 6763 13574
rect 6819 13572 6843 13574
rect 6899 13572 6923 13574
rect 6979 13572 6985 13574
rect 6677 13563 6985 13572
rect 7024 13530 7052 14758
rect 7208 14346 7236 14758
rect 7196 14340 7248 14346
rect 7196 14282 7248 14288
rect 7337 14172 7645 14181
rect 7337 14170 7343 14172
rect 7399 14170 7423 14172
rect 7479 14170 7503 14172
rect 7559 14170 7583 14172
rect 7639 14170 7645 14172
rect 7399 14118 7401 14170
rect 7581 14118 7583 14170
rect 7337 14116 7343 14118
rect 7399 14116 7423 14118
rect 7479 14116 7503 14118
rect 7559 14116 7583 14118
rect 7639 14116 7645 14118
rect 7337 14107 7645 14116
rect 7760 14074 7788 15846
rect 7840 14952 7892 14958
rect 7840 14894 7892 14900
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7196 14000 7248 14006
rect 7196 13942 7248 13948
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 7012 13524 7064 13530
rect 7012 13466 7064 13472
rect 7116 13462 7144 13874
rect 7208 13802 7236 13942
rect 7196 13796 7248 13802
rect 7196 13738 7248 13744
rect 7104 13456 7156 13462
rect 7104 13398 7156 13404
rect 6460 13184 6512 13190
rect 6460 13126 6512 13132
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 6000 12232 6052 12238
rect 6000 12174 6052 12180
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 5816 11280 5868 11286
rect 5816 11222 5868 11228
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 4620 10736 4672 10742
rect 4620 10678 4672 10684
rect 4632 10062 4660 10678
rect 5080 10668 5132 10674
rect 5080 10610 5132 10616
rect 5092 10062 5120 10610
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 4344 9648 4396 9654
rect 4344 9590 4396 9596
rect 4528 9648 4580 9654
rect 4528 9590 4580 9596
rect 4356 9178 4384 9590
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4436 8356 4488 8362
rect 4436 8298 4488 8304
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 4264 7818 4292 8230
rect 4344 7880 4396 7886
rect 4342 7848 4344 7857
rect 4396 7848 4398 7857
rect 4252 7812 4304 7818
rect 4342 7783 4398 7792
rect 4252 7754 4304 7760
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4252 7336 4304 7342
rect 4250 7304 4252 7313
rect 4304 7304 4306 7313
rect 4250 7239 4306 7248
rect 4068 7200 4120 7206
rect 4068 7142 4120 7148
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 3519 6556 3827 6565
rect 3519 6554 3525 6556
rect 3581 6554 3605 6556
rect 3661 6554 3685 6556
rect 3741 6554 3765 6556
rect 3821 6554 3827 6556
rect 3581 6502 3583 6554
rect 3763 6502 3765 6554
rect 3519 6500 3525 6502
rect 3581 6500 3605 6502
rect 3661 6500 3685 6502
rect 3741 6500 3765 6502
rect 3821 6500 3827 6502
rect 3519 6491 3827 6500
rect 3896 6390 3924 6734
rect 3884 6384 3936 6390
rect 3884 6326 3936 6332
rect 3988 6322 4016 6734
rect 4172 6458 4200 6734
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 4160 6248 4212 6254
rect 3436 6174 4108 6202
rect 4264 6236 4292 7239
rect 4212 6208 4292 6236
rect 4160 6190 4212 6196
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 3160 5766 3280 5794
rect 3160 5710 3188 5766
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 3160 5302 3188 5646
rect 2780 5296 2832 5302
rect 2780 5238 2832 5244
rect 3148 5296 3200 5302
rect 3148 5238 3200 5244
rect 2596 5160 2648 5166
rect 2596 5102 2648 5108
rect 2136 4616 2188 4622
rect 2136 4558 2188 4564
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2608 4554 2636 5102
rect 2859 4924 3167 4933
rect 2859 4922 2865 4924
rect 2921 4922 2945 4924
rect 3001 4922 3025 4924
rect 3081 4922 3105 4924
rect 3161 4922 3167 4924
rect 2921 4870 2923 4922
rect 3103 4870 3105 4922
rect 2859 4868 2865 4870
rect 2921 4868 2945 4870
rect 3001 4868 3025 4870
rect 3081 4868 3105 4870
rect 3161 4868 3167 4870
rect 2859 4859 3167 4868
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2596 4548 2648 4554
rect 2596 4490 2648 4496
rect 2792 4214 2820 4626
rect 3332 4480 3384 4486
rect 3332 4422 3384 4428
rect 3344 4214 3372 4422
rect 2780 4208 2832 4214
rect 2780 4150 2832 4156
rect 3332 4208 3384 4214
rect 3332 4150 3384 4156
rect 3344 4026 3372 4150
rect 3252 4010 3372 4026
rect 3240 4004 3372 4010
rect 3292 3998 3372 4004
rect 3240 3946 3292 3952
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 2859 3836 3167 3845
rect 2859 3834 2865 3836
rect 2921 3834 2945 3836
rect 3001 3834 3025 3836
rect 3081 3834 3105 3836
rect 3161 3834 3167 3836
rect 2921 3782 2923 3834
rect 3103 3782 3105 3834
rect 2859 3780 2865 3782
rect 2921 3780 2945 3782
rect 3001 3780 3025 3782
rect 3081 3780 3105 3782
rect 3161 3780 3167 3782
rect 2859 3771 3167 3780
rect 3344 3194 3372 3878
rect 3436 3602 3464 6054
rect 3519 5468 3827 5477
rect 3519 5466 3525 5468
rect 3581 5466 3605 5468
rect 3661 5466 3685 5468
rect 3741 5466 3765 5468
rect 3821 5466 3827 5468
rect 3581 5414 3583 5466
rect 3763 5414 3765 5466
rect 3519 5412 3525 5414
rect 3581 5412 3605 5414
rect 3661 5412 3685 5414
rect 3741 5412 3765 5414
rect 3821 5412 3827 5414
rect 3519 5403 3827 5412
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 3528 4826 3556 5102
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3519 4380 3827 4389
rect 3519 4378 3525 4380
rect 3581 4378 3605 4380
rect 3661 4378 3685 4380
rect 3741 4378 3765 4380
rect 3821 4378 3827 4380
rect 3581 4326 3583 4378
rect 3763 4326 3765 4378
rect 3519 4324 3525 4326
rect 3581 4324 3605 4326
rect 3661 4324 3685 4326
rect 3741 4324 3765 4326
rect 3821 4324 3827 4326
rect 3519 4315 3827 4324
rect 3896 4282 3924 6054
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3988 4826 4016 4966
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 3884 4276 3936 4282
rect 3884 4218 3936 4224
rect 4080 4146 4108 6174
rect 4172 5710 4200 6190
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 4356 5370 4384 7686
rect 4448 7426 4476 8298
rect 4540 8072 4568 9590
rect 5552 8974 5580 10202
rect 5644 10130 5672 10406
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5552 8634 5580 8910
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 4620 8084 4672 8090
rect 4540 8044 4620 8072
rect 4620 8026 4672 8032
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4448 7410 4568 7426
rect 4448 7404 4580 7410
rect 4448 7398 4528 7404
rect 4528 7346 4580 7352
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4448 6202 4476 6734
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4540 6322 4568 6598
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4448 6174 4568 6202
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 4448 5642 4476 6054
rect 4540 5710 4568 6174
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4436 5636 4488 5642
rect 4436 5578 4488 5584
rect 4540 5370 4568 5646
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4528 5364 4580 5370
rect 4528 5306 4580 5312
rect 4252 5228 4304 5234
rect 4252 5170 4304 5176
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 4172 4622 4200 4966
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 4264 4078 4292 5170
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4356 4146 4384 4422
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4252 4072 4304 4078
rect 4252 4014 4304 4020
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 4436 3936 4488 3942
rect 4436 3878 4488 3884
rect 3424 3596 3476 3602
rect 3424 3538 3476 3544
rect 3519 3292 3827 3301
rect 3519 3290 3525 3292
rect 3581 3290 3605 3292
rect 3661 3290 3685 3292
rect 3741 3290 3765 3292
rect 3821 3290 3827 3292
rect 3581 3238 3583 3290
rect 3763 3238 3765 3290
rect 3519 3236 3525 3238
rect 3581 3236 3605 3238
rect 3661 3236 3685 3238
rect 3741 3236 3765 3238
rect 3821 3236 3827 3238
rect 3519 3227 3827 3236
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3988 2990 4016 3878
rect 4448 3602 4476 3878
rect 4436 3596 4488 3602
rect 4436 3538 4488 3544
rect 4632 3466 4660 7890
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 4908 7546 4936 7822
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4724 6866 4752 7142
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4816 6798 4844 7142
rect 4804 6792 4856 6798
rect 4804 6734 4856 6740
rect 4712 6452 4764 6458
rect 4816 6440 4844 6734
rect 4764 6412 4844 6440
rect 4712 6394 4764 6400
rect 4816 5710 4844 6412
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4908 4282 4936 7142
rect 5368 6798 5396 8026
rect 5552 8022 5580 8434
rect 5644 8362 5672 10066
rect 5736 10062 5764 10746
rect 5828 10062 5856 11222
rect 5920 10606 5948 12174
rect 6196 11098 6224 12174
rect 6472 11354 6500 13126
rect 6564 12986 6592 13126
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 7116 12782 7144 13398
rect 7208 13326 7236 13738
rect 7300 13530 7328 14010
rect 7564 13932 7616 13938
rect 7564 13874 7616 13880
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 7576 13530 7604 13874
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7564 13524 7616 13530
rect 7564 13466 7616 13472
rect 7380 13456 7432 13462
rect 7432 13416 7512 13444
rect 7380 13398 7432 13404
rect 7484 13410 7512 13416
rect 7668 13410 7696 13874
rect 7484 13382 7696 13410
rect 7668 13326 7696 13382
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 7656 13320 7708 13326
rect 7656 13262 7708 13268
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 7208 12764 7236 13262
rect 7337 13084 7645 13093
rect 7337 13082 7343 13084
rect 7399 13082 7423 13084
rect 7479 13082 7503 13084
rect 7559 13082 7583 13084
rect 7639 13082 7645 13084
rect 7399 13030 7401 13082
rect 7581 13030 7583 13082
rect 7337 13028 7343 13030
rect 7399 13028 7423 13030
rect 7479 13028 7503 13030
rect 7559 13028 7583 13030
rect 7639 13028 7645 13030
rect 7337 13019 7645 13028
rect 7852 12850 7880 14894
rect 8024 14340 8076 14346
rect 8024 14282 8076 14288
rect 8036 13870 8064 14282
rect 8024 13864 8076 13870
rect 8024 13806 8076 13812
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 8128 12986 8156 13126
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 8220 12866 8248 16118
rect 8852 14476 8904 14482
rect 8852 14418 8904 14424
rect 8864 13870 8892 14418
rect 8956 14074 8984 16526
rect 9876 16454 9904 17070
rect 10140 16788 10192 16794
rect 10140 16730 10192 16736
rect 9864 16448 9916 16454
rect 9864 16390 9916 16396
rect 10152 15978 10180 16730
rect 10336 16674 10364 17138
rect 10428 16794 10456 17138
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 12072 17128 12124 17134
rect 12072 17070 12124 17076
rect 10495 16892 10803 16901
rect 10495 16890 10501 16892
rect 10557 16890 10581 16892
rect 10637 16890 10661 16892
rect 10717 16890 10741 16892
rect 10797 16890 10803 16892
rect 10557 16838 10559 16890
rect 10739 16838 10741 16890
rect 10495 16836 10501 16838
rect 10557 16836 10581 16838
rect 10637 16836 10661 16838
rect 10717 16836 10741 16838
rect 10797 16836 10803 16838
rect 10495 16827 10803 16836
rect 10416 16788 10468 16794
rect 10416 16730 10468 16736
rect 10508 16788 10560 16794
rect 10508 16730 10560 16736
rect 10520 16674 10548 16730
rect 10336 16646 10548 16674
rect 10232 16584 10284 16590
rect 10232 16526 10284 16532
rect 10324 16584 10376 16590
rect 10324 16526 10376 16532
rect 10244 16046 10272 16526
rect 10336 16182 10364 16526
rect 10324 16176 10376 16182
rect 10324 16118 10376 16124
rect 10232 16040 10284 16046
rect 10232 15982 10284 15988
rect 10140 15972 10192 15978
rect 10140 15914 10192 15920
rect 9404 15632 9456 15638
rect 9404 15574 9456 15580
rect 9416 15366 9444 15574
rect 9404 15360 9456 15366
rect 9404 15302 9456 15308
rect 9416 14618 9444 15302
rect 10152 14822 10180 15914
rect 10336 15502 10364 16118
rect 10428 15910 10456 16646
rect 10888 16522 10916 17070
rect 11612 16992 11664 16998
rect 11612 16934 11664 16940
rect 10876 16516 10928 16522
rect 10876 16458 10928 16464
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 11072 16114 11100 16390
rect 11155 16348 11463 16357
rect 11155 16346 11161 16348
rect 11217 16346 11241 16348
rect 11297 16346 11321 16348
rect 11377 16346 11401 16348
rect 11457 16346 11463 16348
rect 11217 16294 11219 16346
rect 11399 16294 11401 16346
rect 11155 16292 11161 16294
rect 11217 16292 11241 16294
rect 11297 16292 11321 16294
rect 11377 16292 11401 16294
rect 11457 16292 11463 16294
rect 11155 16283 11463 16292
rect 11624 16114 11652 16934
rect 12084 16794 12112 17070
rect 12176 16794 12204 17138
rect 12624 17060 12676 17066
rect 12624 17002 12676 17008
rect 12072 16788 12124 16794
rect 12072 16730 12124 16736
rect 12164 16788 12216 16794
rect 12164 16730 12216 16736
rect 11888 16448 11940 16454
rect 11888 16390 11940 16396
rect 11900 16250 11928 16390
rect 11888 16244 11940 16250
rect 11888 16186 11940 16192
rect 12084 16182 12112 16730
rect 12532 16720 12584 16726
rect 12532 16662 12584 16668
rect 12072 16176 12124 16182
rect 12072 16118 12124 16124
rect 12544 16114 12572 16662
rect 12636 16590 12664 17002
rect 12624 16584 12676 16590
rect 12624 16526 12676 16532
rect 12716 16584 12768 16590
rect 12716 16526 12768 16532
rect 12728 16250 12756 16526
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 11612 16108 11664 16114
rect 11612 16050 11664 16056
rect 12532 16108 12584 16114
rect 12532 16050 12584 16056
rect 12820 15978 12848 17138
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12912 16658 12940 16934
rect 14200 16794 14228 17138
rect 14313 16892 14621 16901
rect 14313 16890 14319 16892
rect 14375 16890 14399 16892
rect 14455 16890 14479 16892
rect 14535 16890 14559 16892
rect 14615 16890 14621 16892
rect 14375 16838 14377 16890
rect 14557 16838 14559 16890
rect 14313 16836 14319 16838
rect 14375 16836 14399 16838
rect 14455 16836 14479 16838
rect 14535 16836 14559 16838
rect 14615 16836 14621 16838
rect 14313 16827 14621 16836
rect 15028 16794 15056 17138
rect 14188 16788 14240 16794
rect 14188 16730 14240 16736
rect 15016 16788 15068 16794
rect 15016 16730 15068 16736
rect 12900 16652 12952 16658
rect 12900 16594 12952 16600
rect 14372 16652 14424 16658
rect 14372 16594 14424 16600
rect 13728 16584 13780 16590
rect 13728 16526 13780 16532
rect 12900 16448 12952 16454
rect 12900 16390 12952 16396
rect 13636 16448 13688 16454
rect 13636 16390 13688 16396
rect 12912 16250 12940 16390
rect 13648 16250 13676 16390
rect 12900 16244 12952 16250
rect 12900 16186 12952 16192
rect 13636 16244 13688 16250
rect 13636 16186 13688 16192
rect 12808 15972 12860 15978
rect 12808 15914 12860 15920
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10495 15804 10803 15813
rect 10495 15802 10501 15804
rect 10557 15802 10581 15804
rect 10637 15802 10661 15804
rect 10717 15802 10741 15804
rect 10797 15802 10803 15804
rect 10557 15750 10559 15802
rect 10739 15750 10741 15802
rect 10495 15748 10501 15750
rect 10557 15748 10581 15750
rect 10637 15748 10661 15750
rect 10717 15748 10741 15750
rect 10797 15748 10803 15750
rect 10495 15739 10803 15748
rect 12912 15722 12940 16186
rect 13740 16182 13768 16526
rect 13728 16176 13780 16182
rect 13728 16118 13780 16124
rect 13912 16176 13964 16182
rect 13912 16118 13964 16124
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 12728 15694 12940 15722
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 12728 15366 12756 15694
rect 10232 15360 10284 15366
rect 10232 15302 10284 15308
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 10244 15094 10272 15302
rect 11155 15260 11463 15269
rect 11155 15258 11161 15260
rect 11217 15258 11241 15260
rect 11297 15258 11321 15260
rect 11377 15258 11401 15260
rect 11457 15258 11463 15260
rect 11217 15206 11219 15258
rect 11399 15206 11401 15258
rect 11155 15204 11161 15206
rect 11217 15204 11241 15206
rect 11297 15204 11321 15206
rect 11377 15204 11401 15206
rect 11457 15204 11463 15206
rect 11155 15195 11463 15204
rect 12728 15094 12756 15302
rect 10232 15088 10284 15094
rect 10232 15030 10284 15036
rect 12716 15088 12768 15094
rect 12716 15030 12768 15036
rect 10600 15020 10652 15026
rect 10600 14962 10652 14968
rect 10612 14822 10640 14962
rect 13832 14958 13860 15846
rect 13924 15026 13952 16118
rect 14384 15978 14412 16594
rect 14973 16348 15281 16357
rect 14973 16346 14979 16348
rect 15035 16346 15059 16348
rect 15115 16346 15139 16348
rect 15195 16346 15219 16348
rect 15275 16346 15281 16348
rect 15035 16294 15037 16346
rect 15217 16294 15219 16346
rect 14973 16292 14979 16294
rect 15035 16292 15059 16294
rect 15115 16292 15139 16294
rect 15195 16292 15219 16294
rect 15275 16292 15281 16294
rect 14973 16283 15281 16292
rect 14372 15972 14424 15978
rect 14372 15914 14424 15920
rect 14188 15904 14240 15910
rect 14188 15846 14240 15852
rect 14096 15428 14148 15434
rect 14096 15370 14148 15376
rect 13912 15020 13964 15026
rect 13912 14962 13964 14968
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 10140 14816 10192 14822
rect 10140 14758 10192 14764
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12992 14816 13044 14822
rect 12992 14758 13044 14764
rect 10060 14618 10088 14758
rect 10495 14716 10803 14725
rect 10495 14714 10501 14716
rect 10557 14714 10581 14716
rect 10637 14714 10661 14716
rect 10717 14714 10741 14716
rect 10797 14714 10803 14716
rect 10557 14662 10559 14714
rect 10739 14662 10741 14714
rect 10495 14660 10501 14662
rect 10557 14660 10581 14662
rect 10637 14660 10661 14662
rect 10717 14660 10741 14662
rect 10797 14660 10803 14662
rect 10495 14651 10803 14660
rect 10980 14618 11008 14758
rect 12820 14618 12848 14758
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 9232 14006 9260 14350
rect 9680 14340 9732 14346
rect 9680 14282 9732 14288
rect 10600 14340 10652 14346
rect 10600 14282 10652 14288
rect 10784 14340 10836 14346
rect 10784 14282 10836 14288
rect 10876 14340 10928 14346
rect 10876 14282 10928 14288
rect 9692 14074 9720 14282
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9784 14074 9812 14214
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9220 14000 9272 14006
rect 9220 13942 9272 13948
rect 10612 13938 10640 14282
rect 9128 13932 9180 13938
rect 9128 13874 9180 13880
rect 10600 13932 10652 13938
rect 10796 13920 10824 14282
rect 10888 14074 10916 14282
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 10876 13932 10928 13938
rect 10796 13892 10876 13920
rect 10600 13874 10652 13880
rect 10876 13874 10928 13880
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 8576 13864 8628 13870
rect 8576 13806 8628 13812
rect 8852 13864 8904 13870
rect 8852 13806 8904 13812
rect 8404 13530 8432 13806
rect 8588 13530 8616 13806
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 8404 13326 8432 13466
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 8300 13252 8352 13258
rect 8300 13194 8352 13200
rect 8312 12986 8340 13194
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8220 12850 8340 12866
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7840 12844 7892 12850
rect 7840 12786 7892 12792
rect 7932 12844 7984 12850
rect 8220 12844 8352 12850
rect 8220 12838 8300 12844
rect 7984 12804 8064 12832
rect 7932 12786 7984 12792
rect 7288 12776 7340 12782
rect 7208 12736 7288 12764
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6564 12434 6592 12582
rect 6677 12540 6985 12549
rect 6677 12538 6683 12540
rect 6739 12538 6763 12540
rect 6819 12538 6843 12540
rect 6899 12538 6923 12540
rect 6979 12538 6985 12540
rect 6739 12486 6741 12538
rect 6921 12486 6923 12538
rect 6677 12484 6683 12486
rect 6739 12484 6763 12486
rect 6819 12484 6843 12486
rect 6899 12484 6923 12486
rect 6979 12484 6985 12486
rect 6677 12475 6985 12484
rect 6564 12406 6684 12434
rect 6552 12164 6604 12170
rect 6552 12106 6604 12112
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6104 11070 6224 11098
rect 6104 10810 6132 11070
rect 6184 11008 6236 11014
rect 6184 10950 6236 10956
rect 6276 11008 6328 11014
rect 6276 10950 6328 10956
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6092 10804 6144 10810
rect 6092 10746 6144 10752
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 6092 10668 6144 10674
rect 6092 10610 6144 10616
rect 5908 10600 5960 10606
rect 5908 10542 5960 10548
rect 6012 10266 6040 10610
rect 6104 10266 6132 10610
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 5908 10192 5960 10198
rect 6196 10146 6224 10950
rect 6288 10606 6316 10950
rect 6368 10736 6420 10742
rect 6368 10678 6420 10684
rect 6276 10600 6328 10606
rect 6276 10542 6328 10548
rect 5908 10134 5960 10140
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5920 9926 5948 10134
rect 6104 10118 6224 10146
rect 6380 10130 6408 10678
rect 6368 10124 6420 10130
rect 6104 10062 6132 10118
rect 6368 10066 6420 10072
rect 6472 10062 6500 10950
rect 6564 10674 6592 12106
rect 6656 11558 6684 12406
rect 7104 12368 7156 12374
rect 7104 12310 7156 12316
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6677 11452 6985 11461
rect 6677 11450 6683 11452
rect 6739 11450 6763 11452
rect 6819 11450 6843 11452
rect 6899 11450 6923 11452
rect 6979 11450 6985 11452
rect 6739 11398 6741 11450
rect 6921 11398 6923 11450
rect 6677 11396 6683 11398
rect 6739 11396 6763 11398
rect 6819 11396 6843 11398
rect 6899 11396 6923 11398
rect 6979 11396 6985 11398
rect 6677 11387 6985 11396
rect 7116 11354 7144 12310
rect 7208 11830 7236 12736
rect 7288 12718 7340 12724
rect 7484 12238 7512 12786
rect 7852 12646 7880 12786
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7337 11996 7645 12005
rect 7337 11994 7343 11996
rect 7399 11994 7423 11996
rect 7479 11994 7503 11996
rect 7559 11994 7583 11996
rect 7639 11994 7645 11996
rect 7399 11942 7401 11994
rect 7581 11942 7583 11994
rect 7337 11940 7343 11942
rect 7399 11940 7423 11942
rect 7479 11940 7503 11942
rect 7559 11940 7583 11942
rect 7639 11940 7645 11942
rect 7337 11931 7645 11940
rect 7196 11824 7248 11830
rect 7196 11766 7248 11772
rect 7564 11824 7616 11830
rect 7564 11766 7616 11772
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6748 10452 6776 11154
rect 7116 11082 7144 11290
rect 7484 11150 7512 11494
rect 7576 11150 7604 11766
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7668 11150 7696 11494
rect 7760 11286 7788 12242
rect 7852 12238 7880 12582
rect 8036 12374 8064 12804
rect 8300 12786 8352 12792
rect 8312 12714 8340 12786
rect 8300 12708 8352 12714
rect 8300 12650 8352 12656
rect 8024 12368 8076 12374
rect 8024 12310 8076 12316
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7564 11144 7616 11150
rect 7564 11086 7616 11092
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7104 11076 7156 11082
rect 7104 11018 7156 11024
rect 7484 11014 7512 11086
rect 7760 11082 7788 11222
rect 7748 11076 7800 11082
rect 7748 11018 7800 11024
rect 7472 11008 7524 11014
rect 7472 10950 7524 10956
rect 7337 10908 7645 10917
rect 7337 10906 7343 10908
rect 7399 10906 7423 10908
rect 7479 10906 7503 10908
rect 7559 10906 7583 10908
rect 7639 10906 7645 10908
rect 7399 10854 7401 10906
rect 7581 10854 7583 10906
rect 7337 10852 7343 10854
rect 7399 10852 7423 10854
rect 7479 10852 7503 10854
rect 7559 10852 7583 10854
rect 7639 10852 7645 10854
rect 7337 10843 7645 10852
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 6564 10424 6776 10452
rect 6564 10062 6592 10424
rect 6677 10364 6985 10373
rect 6677 10362 6683 10364
rect 6739 10362 6763 10364
rect 6819 10362 6843 10364
rect 6899 10362 6923 10364
rect 6979 10362 6985 10364
rect 6739 10310 6741 10362
rect 6921 10310 6923 10362
rect 6677 10308 6683 10310
rect 6739 10308 6763 10310
rect 6819 10308 6843 10310
rect 6899 10308 6923 10310
rect 6979 10308 6985 10310
rect 6677 10299 6985 10308
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 5908 9920 5960 9926
rect 5908 9862 5960 9868
rect 5908 9104 5960 9110
rect 5908 9046 5960 9052
rect 5724 8900 5776 8906
rect 5724 8842 5776 8848
rect 5736 8498 5764 8842
rect 5920 8498 5948 9046
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 6012 8498 6040 8842
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 5540 8016 5592 8022
rect 5540 7958 5592 7964
rect 5552 7546 5580 7958
rect 6012 7698 6040 8434
rect 5828 7670 6040 7698
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5828 7410 5856 7670
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5460 7313 5488 7346
rect 5446 7304 5502 7313
rect 5502 7262 5580 7290
rect 5446 7239 5502 7248
rect 5552 6934 5580 7262
rect 5828 7206 5856 7346
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5540 6928 5592 6934
rect 5540 6870 5592 6876
rect 5552 6798 5580 6870
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 4988 6384 5040 6390
rect 4988 6326 5040 6332
rect 5000 5914 5028 6326
rect 4988 5908 5040 5914
rect 4988 5850 5040 5856
rect 5092 5234 5120 6598
rect 5276 6254 5304 6598
rect 5368 6254 5396 6734
rect 5644 6730 5672 7142
rect 5828 7002 5856 7142
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 5632 6724 5684 6730
rect 5632 6666 5684 6672
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5644 5846 5672 6666
rect 5920 6322 5948 7482
rect 6104 7002 6132 9998
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6196 8498 6224 8978
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 6472 7546 6500 9318
rect 6564 9110 6592 9998
rect 6932 9654 6960 9998
rect 7012 9716 7064 9722
rect 7012 9658 7064 9664
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 6677 9276 6985 9285
rect 6677 9274 6683 9276
rect 6739 9274 6763 9276
rect 6819 9274 6843 9276
rect 6899 9274 6923 9276
rect 6979 9274 6985 9276
rect 6739 9222 6741 9274
rect 6921 9222 6923 9274
rect 6677 9220 6683 9222
rect 6739 9220 6763 9222
rect 6819 9220 6843 9222
rect 6899 9220 6923 9222
rect 6979 9220 6985 9222
rect 6677 9211 6985 9220
rect 6552 9104 6604 9110
rect 6552 9046 6604 9052
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6564 8566 6592 8910
rect 6748 8634 6776 8910
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6552 8560 6604 8566
rect 6552 8502 6604 8508
rect 7024 8430 7052 9658
rect 7012 8424 7064 8430
rect 7012 8366 7064 8372
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 6677 8188 6985 8197
rect 6677 8186 6683 8188
rect 6739 8186 6763 8188
rect 6819 8186 6843 8188
rect 6899 8186 6923 8188
rect 6979 8186 6985 8188
rect 6739 8134 6741 8186
rect 6921 8134 6923 8186
rect 6677 8132 6683 8134
rect 6739 8132 6763 8134
rect 6819 8132 6843 8134
rect 6899 8132 6923 8134
rect 6979 8132 6985 8134
rect 6677 8123 6985 8132
rect 7024 7886 7052 8230
rect 6828 7880 6880 7886
rect 7012 7880 7064 7886
rect 6880 7840 7012 7868
rect 6828 7822 6880 7828
rect 7012 7822 7064 7828
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 7024 7274 7052 7822
rect 7012 7268 7064 7274
rect 7012 7210 7064 7216
rect 6184 7200 6236 7206
rect 6184 7142 6236 7148
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6196 7002 6224 7142
rect 6092 6996 6144 7002
rect 6092 6938 6144 6944
rect 6184 6996 6236 7002
rect 6184 6938 6236 6944
rect 6460 6928 6512 6934
rect 6460 6870 6512 6876
rect 6368 6860 6420 6866
rect 6368 6802 6420 6808
rect 6380 6322 6408 6802
rect 6472 6322 6500 6870
rect 6564 6440 6592 7142
rect 6677 7100 6985 7109
rect 6677 7098 6683 7100
rect 6739 7098 6763 7100
rect 6819 7098 6843 7100
rect 6899 7098 6923 7100
rect 6979 7098 6985 7100
rect 6739 7046 6741 7098
rect 6921 7046 6923 7098
rect 6677 7044 6683 7046
rect 6739 7044 6763 7046
rect 6819 7044 6843 7046
rect 6899 7044 6923 7046
rect 6979 7044 6985 7046
rect 6677 7035 6985 7044
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6828 6724 6880 6730
rect 6828 6666 6880 6672
rect 6564 6412 6776 6440
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6000 6180 6052 6186
rect 6000 6122 6052 6128
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5632 5840 5684 5846
rect 5632 5782 5684 5788
rect 5828 5778 5856 6054
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 6012 5710 6040 6122
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6104 5710 6132 5850
rect 6196 5710 6224 6258
rect 6564 5914 6592 6412
rect 6748 6322 6776 6412
rect 6840 6390 6868 6666
rect 6828 6384 6880 6390
rect 6828 6326 6880 6332
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6656 6186 6684 6258
rect 6644 6180 6696 6186
rect 6644 6122 6696 6128
rect 6932 6100 6960 6802
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 7024 6458 7052 6598
rect 7116 6458 7144 10542
rect 7760 10470 7788 11018
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 7337 9820 7645 9829
rect 7337 9818 7343 9820
rect 7399 9818 7423 9820
rect 7479 9818 7503 9820
rect 7559 9818 7583 9820
rect 7639 9818 7645 9820
rect 7399 9766 7401 9818
rect 7581 9766 7583 9818
rect 7337 9764 7343 9766
rect 7399 9764 7423 9766
rect 7479 9764 7503 9766
rect 7559 9764 7583 9766
rect 7639 9764 7645 9766
rect 7337 9755 7645 9764
rect 7852 9674 7880 12174
rect 7932 11008 7984 11014
rect 7932 10950 7984 10956
rect 7564 9648 7616 9654
rect 7470 9616 7526 9625
rect 7392 9586 7470 9602
rect 7380 9580 7470 9586
rect 7432 9574 7470 9580
rect 7564 9590 7616 9596
rect 7668 9646 7880 9674
rect 7470 9551 7526 9560
rect 7380 9522 7432 9528
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 7208 8362 7236 9454
rect 7472 9444 7524 9450
rect 7472 9386 7524 9392
rect 7484 9110 7512 9386
rect 7472 9104 7524 9110
rect 7470 9072 7472 9081
rect 7524 9072 7526 9081
rect 7470 9007 7526 9016
rect 7576 8974 7604 9590
rect 7668 9586 7696 9646
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7668 9042 7696 9522
rect 7656 9036 7708 9042
rect 7708 8996 7788 9024
rect 7656 8978 7708 8984
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 7337 8732 7645 8741
rect 7337 8730 7343 8732
rect 7399 8730 7423 8732
rect 7479 8730 7503 8732
rect 7559 8730 7583 8732
rect 7639 8730 7645 8732
rect 7399 8678 7401 8730
rect 7581 8678 7583 8730
rect 7337 8676 7343 8678
rect 7399 8676 7423 8678
rect 7479 8676 7503 8678
rect 7559 8676 7583 8678
rect 7639 8676 7645 8678
rect 7337 8667 7645 8676
rect 7760 8634 7788 8996
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 7196 8356 7248 8362
rect 7196 8298 7248 8304
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 6932 6072 7052 6100
rect 6677 6012 6985 6021
rect 6677 6010 6683 6012
rect 6739 6010 6763 6012
rect 6819 6010 6843 6012
rect 6899 6010 6923 6012
rect 6979 6010 6985 6012
rect 6739 5958 6741 6010
rect 6921 5958 6923 6010
rect 6677 5956 6683 5958
rect 6739 5956 6763 5958
rect 6819 5956 6843 5958
rect 6899 5956 6923 5958
rect 6979 5956 6985 5958
rect 6677 5947 6985 5956
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 6368 5772 6420 5778
rect 6368 5714 6420 5720
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6012 5574 6040 5646
rect 6000 5568 6052 5574
rect 6000 5510 6052 5516
rect 6380 5234 6408 5714
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 5368 3738 5396 5102
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 6104 4758 6132 4966
rect 6380 4758 6408 5170
rect 6677 4924 6985 4933
rect 6677 4922 6683 4924
rect 6739 4922 6763 4924
rect 6819 4922 6843 4924
rect 6899 4922 6923 4924
rect 6979 4922 6985 4924
rect 6739 4870 6741 4922
rect 6921 4870 6923 4922
rect 6677 4868 6683 4870
rect 6739 4868 6763 4870
rect 6819 4868 6843 4870
rect 6899 4868 6923 4870
rect 6979 4868 6985 4870
rect 6677 4859 6985 4868
rect 7024 4826 7052 6072
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 6092 4752 6144 4758
rect 6092 4694 6144 4700
rect 6368 4752 6420 4758
rect 6368 4694 6420 4700
rect 7104 4616 7156 4622
rect 7024 4576 7104 4604
rect 7024 4146 7052 4576
rect 7104 4558 7156 4564
rect 7208 4434 7236 7822
rect 7300 7818 7328 8366
rect 7484 7886 7512 8434
rect 7852 8090 7880 8774
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7288 7812 7340 7818
rect 7288 7754 7340 7760
rect 7337 7644 7645 7653
rect 7337 7642 7343 7644
rect 7399 7642 7423 7644
rect 7479 7642 7503 7644
rect 7559 7642 7583 7644
rect 7639 7642 7645 7644
rect 7399 7590 7401 7642
rect 7581 7590 7583 7642
rect 7337 7588 7343 7590
rect 7399 7588 7423 7590
rect 7479 7588 7503 7590
rect 7559 7588 7583 7590
rect 7639 7588 7645 7590
rect 7337 7579 7645 7588
rect 7564 7540 7616 7546
rect 7944 7528 7972 10950
rect 8036 9382 8064 12174
rect 8312 11642 8340 12650
rect 8404 12442 8432 13262
rect 8864 12986 8892 13806
rect 9140 13530 9168 13874
rect 10495 13628 10803 13637
rect 10495 13626 10501 13628
rect 10557 13626 10581 13628
rect 10637 13626 10661 13628
rect 10717 13626 10741 13628
rect 10797 13626 10803 13628
rect 10557 13574 10559 13626
rect 10739 13574 10741 13626
rect 10495 13572 10501 13574
rect 10557 13572 10581 13574
rect 10637 13572 10661 13574
rect 10717 13572 10741 13574
rect 10797 13572 10803 13574
rect 10495 13563 10803 13572
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 10888 13326 10916 13874
rect 11072 13462 11100 14214
rect 11155 14172 11463 14181
rect 11155 14170 11161 14172
rect 11217 14170 11241 14172
rect 11297 14170 11321 14172
rect 11377 14170 11401 14172
rect 11457 14170 11463 14172
rect 11217 14118 11219 14170
rect 11399 14118 11401 14170
rect 11155 14116 11161 14118
rect 11217 14116 11241 14118
rect 11297 14116 11321 14118
rect 11377 14116 11401 14118
rect 11457 14116 11463 14118
rect 11155 14107 11463 14116
rect 12348 13524 12400 13530
rect 12348 13466 12400 13472
rect 11060 13456 11112 13462
rect 11060 13398 11112 13404
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 11520 13320 11572 13326
rect 11520 13262 11572 13268
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 10152 12986 10180 13262
rect 10324 13252 10376 13258
rect 10324 13194 10376 13200
rect 8852 12980 8904 12986
rect 8852 12922 8904 12928
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 9128 12912 9180 12918
rect 9128 12854 9180 12860
rect 8576 12640 8628 12646
rect 8576 12582 8628 12588
rect 8392 12436 8444 12442
rect 8392 12378 8444 12384
rect 8484 11688 8536 11694
rect 8312 11614 8432 11642
rect 8484 11630 8536 11636
rect 8404 10470 8432 11614
rect 8496 11150 8524 11630
rect 8588 11558 8616 12582
rect 9036 12300 9088 12306
rect 9036 12242 9088 12248
rect 9048 11898 9076 12242
rect 9140 12238 9168 12854
rect 10336 12850 10364 13194
rect 10704 12986 10732 13262
rect 11155 13084 11463 13093
rect 11155 13082 11161 13084
rect 11217 13082 11241 13084
rect 11297 13082 11321 13084
rect 11377 13082 11401 13084
rect 11457 13082 11463 13084
rect 11217 13030 11219 13082
rect 11399 13030 11401 13082
rect 11155 13028 11161 13030
rect 11217 13028 11241 13030
rect 11297 13028 11321 13030
rect 11377 13028 11401 13030
rect 11457 13028 11463 13030
rect 11155 13019 11463 13028
rect 11532 12986 11560 13262
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 10324 12844 10376 12850
rect 10324 12786 10376 12792
rect 11624 12782 11652 13262
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 11612 12776 11664 12782
rect 11612 12718 11664 12724
rect 10060 12442 10088 12718
rect 12072 12640 12124 12646
rect 12072 12582 12124 12588
rect 10495 12540 10803 12549
rect 10495 12538 10501 12540
rect 10557 12538 10581 12540
rect 10637 12538 10661 12540
rect 10717 12538 10741 12540
rect 10797 12538 10803 12540
rect 10557 12486 10559 12538
rect 10739 12486 10741 12538
rect 10495 12484 10501 12486
rect 10557 12484 10581 12486
rect 10637 12484 10661 12486
rect 10717 12484 10741 12486
rect 10797 12484 10803 12486
rect 10495 12475 10803 12484
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 11980 12368 12032 12374
rect 11980 12310 12032 12316
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9956 12096 10008 12102
rect 9956 12038 10008 12044
rect 10876 12096 10928 12102
rect 10876 12038 10928 12044
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 8852 11824 8904 11830
rect 8852 11766 8904 11772
rect 8576 11552 8628 11558
rect 8576 11494 8628 11500
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8680 11354 8708 11494
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8864 11150 8892 11766
rect 9968 11762 9996 12038
rect 10888 11898 10916 12038
rect 11155 11996 11463 12005
rect 11155 11994 11161 11996
rect 11217 11994 11241 11996
rect 11297 11994 11321 11996
rect 11377 11994 11401 11996
rect 11457 11994 11463 11996
rect 11217 11942 11219 11994
rect 11399 11942 11401 11994
rect 11155 11940 11161 11942
rect 11217 11940 11241 11942
rect 11297 11940 11321 11942
rect 11377 11940 11401 11942
rect 11457 11940 11463 11942
rect 11155 11931 11463 11940
rect 11992 11898 12020 12310
rect 12084 12238 12112 12582
rect 12360 12442 12388 13466
rect 12728 13326 12756 14214
rect 13004 13530 13032 14758
rect 13924 13530 13952 14962
rect 14108 14958 14136 15370
rect 14200 15366 14228 15846
rect 14313 15804 14621 15813
rect 14313 15802 14319 15804
rect 14375 15802 14399 15804
rect 14455 15802 14479 15804
rect 14535 15802 14559 15804
rect 14615 15802 14621 15804
rect 14375 15750 14377 15802
rect 14557 15750 14559 15802
rect 14313 15748 14319 15750
rect 14375 15748 14399 15750
rect 14455 15748 14479 15750
rect 14535 15748 14559 15750
rect 14615 15748 14621 15750
rect 14313 15739 14621 15748
rect 14188 15360 14240 15366
rect 14188 15302 14240 15308
rect 16028 15360 16080 15366
rect 16028 15302 16080 15308
rect 14200 15026 14228 15302
rect 14973 15260 15281 15269
rect 14973 15258 14979 15260
rect 15035 15258 15059 15260
rect 15115 15258 15139 15260
rect 15195 15258 15219 15260
rect 15275 15258 15281 15260
rect 15035 15206 15037 15258
rect 15217 15206 15219 15258
rect 14973 15204 14979 15206
rect 15035 15204 15059 15206
rect 15115 15204 15139 15206
rect 15195 15204 15219 15206
rect 15275 15204 15281 15206
rect 14973 15195 15281 15204
rect 16040 15065 16068 15302
rect 16026 15056 16082 15065
rect 14188 15020 14240 15026
rect 16026 14991 16082 15000
rect 14188 14962 14240 14968
rect 14096 14952 14148 14958
rect 14096 14894 14148 14900
rect 14313 14716 14621 14725
rect 14313 14714 14319 14716
rect 14375 14714 14399 14716
rect 14455 14714 14479 14716
rect 14535 14714 14559 14716
rect 14615 14714 14621 14716
rect 14375 14662 14377 14714
rect 14557 14662 14559 14714
rect 14313 14660 14319 14662
rect 14375 14660 14399 14662
rect 14455 14660 14479 14662
rect 14535 14660 14559 14662
rect 14615 14660 14621 14662
rect 14313 14651 14621 14660
rect 14973 14172 15281 14181
rect 14973 14170 14979 14172
rect 15035 14170 15059 14172
rect 15115 14170 15139 14172
rect 15195 14170 15219 14172
rect 15275 14170 15281 14172
rect 15035 14118 15037 14170
rect 15217 14118 15219 14170
rect 14973 14116 14979 14118
rect 15035 14116 15059 14118
rect 15115 14116 15139 14118
rect 15195 14116 15219 14118
rect 15275 14116 15281 14118
rect 14973 14107 15281 14116
rect 14313 13628 14621 13637
rect 14313 13626 14319 13628
rect 14375 13626 14399 13628
rect 14455 13626 14479 13628
rect 14535 13626 14559 13628
rect 14615 13626 14621 13628
rect 14375 13574 14377 13626
rect 14557 13574 14559 13626
rect 14313 13572 14319 13574
rect 14375 13572 14399 13574
rect 14455 13572 14479 13574
rect 14535 13572 14559 13574
rect 14615 13572 14621 13574
rect 14313 13563 14621 13572
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 13912 13320 13964 13326
rect 13912 13262 13964 13268
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13648 12850 13676 13126
rect 13636 12844 13688 12850
rect 13636 12786 13688 12792
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 12348 12436 12400 12442
rect 13372 12434 13400 12718
rect 13372 12406 13492 12434
rect 12348 12378 12400 12384
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 13464 12170 13492 12406
rect 13648 12374 13676 12786
rect 13924 12442 13952 13262
rect 14372 13184 14424 13190
rect 14372 13126 14424 13132
rect 14832 13184 14884 13190
rect 14832 13126 14884 13132
rect 14384 12782 14412 13126
rect 14844 12850 14872 13126
rect 14973 13084 15281 13093
rect 14973 13082 14979 13084
rect 15035 13082 15059 13084
rect 15115 13082 15139 13084
rect 15195 13082 15219 13084
rect 15275 13082 15281 13084
rect 15035 13030 15037 13082
rect 15217 13030 15219 13082
rect 14973 13028 14979 13030
rect 15035 13028 15059 13030
rect 15115 13028 15139 13030
rect 15195 13028 15219 13030
rect 15275 13028 15281 13030
rect 14973 13019 15281 13028
rect 15764 12986 15792 13262
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 15948 13025 15976 13126
rect 15934 13016 15990 13025
rect 15752 12980 15804 12986
rect 15934 12951 15990 12960
rect 15752 12922 15804 12928
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 14372 12776 14424 12782
rect 14372 12718 14424 12724
rect 14313 12540 14621 12549
rect 14313 12538 14319 12540
rect 14375 12538 14399 12540
rect 14455 12538 14479 12540
rect 14535 12538 14559 12540
rect 14615 12538 14621 12540
rect 14375 12486 14377 12538
rect 14557 12486 14559 12538
rect 14313 12484 14319 12486
rect 14375 12484 14399 12486
rect 14455 12484 14479 12486
rect 14535 12484 14559 12486
rect 14615 12484 14621 12486
rect 14313 12475 14621 12484
rect 13912 12436 13964 12442
rect 13912 12378 13964 12384
rect 13636 12368 13688 12374
rect 13636 12310 13688 12316
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12912 11898 12940 12038
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 11704 11756 11756 11762
rect 11704 11698 11756 11704
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9692 11286 9720 11562
rect 10495 11452 10803 11461
rect 10495 11450 10501 11452
rect 10557 11450 10581 11452
rect 10637 11450 10661 11452
rect 10717 11450 10741 11452
rect 10797 11450 10803 11452
rect 10557 11398 10559 11450
rect 10739 11398 10741 11450
rect 10495 11396 10501 11398
rect 10557 11396 10581 11398
rect 10637 11396 10661 11398
rect 10717 11396 10741 11398
rect 10797 11396 10803 11398
rect 10495 11387 10803 11396
rect 9680 11280 9732 11286
rect 9680 11222 9732 11228
rect 11532 11150 11560 11698
rect 11716 11286 11744 11698
rect 11704 11280 11756 11286
rect 11704 11222 11756 11228
rect 12268 11150 12296 11834
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8116 9988 8168 9994
rect 8116 9930 8168 9936
rect 8128 9654 8156 9930
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 8220 9722 8248 9862
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 8116 9648 8168 9654
rect 8312 9602 8340 10406
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8404 9654 8432 10202
rect 8576 9988 8628 9994
rect 8576 9930 8628 9936
rect 8588 9654 8616 9930
rect 8116 9590 8168 9596
rect 8220 9574 8340 9602
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 8576 9648 8628 9654
rect 8576 9590 8628 9596
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 8036 8634 8064 9318
rect 8116 9036 8168 9042
rect 8116 8978 8168 8984
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 8128 8090 8156 8978
rect 8220 8566 8248 9574
rect 8392 9104 8444 9110
rect 8390 9072 8392 9081
rect 8444 9072 8446 9081
rect 8390 9007 8446 9016
rect 8588 8974 8616 9590
rect 8864 9058 8892 11086
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9324 10062 9352 10406
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9508 10062 9536 10202
rect 9692 10198 9720 10950
rect 11155 10908 11463 10917
rect 11155 10906 11161 10908
rect 11217 10906 11241 10908
rect 11297 10906 11321 10908
rect 11377 10906 11401 10908
rect 11457 10906 11463 10908
rect 11217 10854 11219 10906
rect 11399 10854 11401 10906
rect 11155 10852 11161 10854
rect 11217 10852 11241 10854
rect 11297 10852 11321 10854
rect 11377 10852 11401 10854
rect 11457 10852 11463 10854
rect 11155 10843 11463 10852
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 9968 10198 9996 10746
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 10495 10364 10803 10373
rect 10495 10362 10501 10364
rect 10557 10362 10581 10364
rect 10637 10362 10661 10364
rect 10717 10362 10741 10364
rect 10797 10362 10803 10364
rect 10557 10310 10559 10362
rect 10739 10310 10741 10362
rect 10495 10308 10501 10310
rect 10557 10308 10581 10310
rect 10637 10308 10661 10310
rect 10717 10308 10741 10310
rect 10797 10308 10803 10310
rect 10495 10299 10803 10308
rect 12360 10266 12388 10542
rect 12728 10266 12756 10610
rect 13372 10606 13400 11086
rect 13464 10810 13492 12106
rect 14844 11898 14872 12786
rect 14973 11996 15281 12005
rect 14973 11994 14979 11996
rect 15035 11994 15059 11996
rect 15115 11994 15139 11996
rect 15195 11994 15219 11996
rect 15275 11994 15281 11996
rect 15035 11942 15037 11994
rect 15217 11942 15219 11994
rect 14973 11940 14979 11942
rect 15035 11940 15059 11942
rect 15115 11940 15139 11942
rect 15195 11940 15219 11942
rect 15275 11940 15281 11942
rect 14973 11931 15281 11940
rect 14832 11892 14884 11898
rect 14832 11834 14884 11840
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 15016 11756 15068 11762
rect 15016 11698 15068 11704
rect 13820 11280 13872 11286
rect 13820 11222 13872 11228
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 13556 10742 13584 11154
rect 13544 10736 13596 10742
rect 13544 10678 13596 10684
rect 13360 10600 13412 10606
rect 13360 10542 13412 10548
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 9680 10192 9732 10198
rect 9680 10134 9732 10140
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9956 10056 10008 10062
rect 9956 9998 10008 10004
rect 12072 10056 12124 10062
rect 12124 10004 12296 10010
rect 12072 9998 12296 10004
rect 9048 9654 9076 9998
rect 9036 9648 9088 9654
rect 9034 9616 9036 9625
rect 9088 9616 9090 9625
rect 9034 9551 9090 9560
rect 9128 9580 9180 9586
rect 8772 9030 8892 9058
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 8116 8084 8168 8090
rect 8116 8026 8168 8032
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 7616 7500 7972 7528
rect 7564 7482 7616 7488
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 7300 7206 7328 7346
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 7576 6934 7604 7346
rect 7840 7268 7892 7274
rect 7840 7210 7892 7216
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7564 6928 7616 6934
rect 7564 6870 7616 6876
rect 7337 6556 7645 6565
rect 7337 6554 7343 6556
rect 7399 6554 7423 6556
rect 7479 6554 7503 6556
rect 7559 6554 7583 6556
rect 7639 6554 7645 6556
rect 7399 6502 7401 6554
rect 7581 6502 7583 6554
rect 7337 6500 7343 6502
rect 7399 6500 7423 6502
rect 7479 6500 7503 6502
rect 7559 6500 7583 6502
rect 7639 6500 7645 6502
rect 7337 6491 7645 6500
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7484 5914 7512 6190
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 7668 5710 7696 6054
rect 7656 5704 7708 5710
rect 7656 5646 7708 5652
rect 7337 5468 7645 5477
rect 7337 5466 7343 5468
rect 7399 5466 7423 5468
rect 7479 5466 7503 5468
rect 7559 5466 7583 5468
rect 7639 5466 7645 5468
rect 7399 5414 7401 5466
rect 7581 5414 7583 5466
rect 7337 5412 7343 5414
rect 7399 5412 7423 5414
rect 7479 5412 7503 5414
rect 7559 5412 7583 5414
rect 7639 5412 7645 5414
rect 7337 5403 7645 5412
rect 7656 4684 7708 4690
rect 7656 4626 7708 4632
rect 7564 4616 7616 4622
rect 7564 4558 7616 4564
rect 7576 4486 7604 4558
rect 7116 4406 7236 4434
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 7668 4434 7696 4626
rect 7668 4406 7701 4434
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 6677 3836 6985 3845
rect 6677 3834 6683 3836
rect 6739 3834 6763 3836
rect 6819 3834 6843 3836
rect 6899 3834 6923 3836
rect 6979 3834 6985 3836
rect 6739 3782 6741 3834
rect 6921 3782 6923 3834
rect 6677 3780 6683 3782
rect 6739 3780 6763 3782
rect 6819 3780 6843 3782
rect 6899 3780 6923 3782
rect 6979 3780 6985 3782
rect 6677 3771 6985 3780
rect 7024 3738 7052 4082
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 4620 3460 4672 3466
rect 4620 3402 4672 3408
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 4172 3194 4200 3334
rect 4632 3194 4660 3402
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 5368 3058 5396 3674
rect 6090 3632 6146 3641
rect 6090 3567 6092 3576
rect 6144 3567 6146 3576
rect 6092 3538 6144 3544
rect 6288 3534 6316 3674
rect 6736 3664 6788 3670
rect 6734 3632 6736 3641
rect 6920 3664 6972 3670
rect 6788 3632 6790 3641
rect 6920 3606 6972 3612
rect 6734 3567 6790 3576
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 6368 3460 6420 3466
rect 6552 3460 6604 3466
rect 6420 3420 6552 3448
rect 6368 3402 6420 3408
rect 6552 3402 6604 3408
rect 5632 3392 5684 3398
rect 5632 3334 5684 3340
rect 5816 3392 5868 3398
rect 5816 3334 5868 3340
rect 5644 3194 5672 3334
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5828 3058 5856 3334
rect 6932 3058 6960 3606
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 7024 3194 7052 3334
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 1952 2984 2004 2990
rect 1952 2926 2004 2932
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 4344 2916 4396 2922
rect 4344 2858 4396 2864
rect 938 2816 994 2825
rect 938 2751 994 2760
rect 2859 2748 3167 2757
rect 2859 2746 2865 2748
rect 2921 2746 2945 2748
rect 3001 2746 3025 2748
rect 3081 2746 3105 2748
rect 3161 2746 3167 2748
rect 2921 2694 2923 2746
rect 3103 2694 3105 2746
rect 2859 2692 2865 2694
rect 2921 2692 2945 2694
rect 3001 2692 3025 2694
rect 3081 2692 3105 2694
rect 3161 2692 3167 2694
rect 2859 2683 3167 2692
rect 4356 2446 4384 2858
rect 6677 2748 6985 2757
rect 6677 2746 6683 2748
rect 6739 2746 6763 2748
rect 6819 2746 6843 2748
rect 6899 2746 6923 2748
rect 6979 2746 6985 2748
rect 6739 2694 6741 2746
rect 6921 2694 6923 2746
rect 6677 2692 6683 2694
rect 6739 2692 6763 2694
rect 6819 2692 6843 2694
rect 6899 2692 6923 2694
rect 6979 2692 6985 2694
rect 6677 2683 6985 2692
rect 7116 2650 7144 4406
rect 7337 4380 7645 4389
rect 7337 4378 7343 4380
rect 7399 4378 7423 4380
rect 7479 4378 7503 4380
rect 7559 4378 7583 4380
rect 7639 4378 7645 4380
rect 7399 4326 7401 4378
rect 7581 4326 7583 4378
rect 7337 4324 7343 4326
rect 7399 4324 7423 4326
rect 7479 4324 7503 4326
rect 7559 4324 7583 4326
rect 7639 4324 7645 4326
rect 7337 4315 7645 4324
rect 7673 4298 7701 4406
rect 7668 4270 7701 4298
rect 7668 4078 7696 4270
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7208 2990 7236 3878
rect 7337 3292 7645 3301
rect 7337 3290 7343 3292
rect 7399 3290 7423 3292
rect 7479 3290 7503 3292
rect 7559 3290 7583 3292
rect 7639 3290 7645 3292
rect 7399 3238 7401 3290
rect 7581 3238 7583 3290
rect 7337 3236 7343 3238
rect 7399 3236 7423 3238
rect 7479 3236 7503 3238
rect 7559 3236 7583 3238
rect 7639 3236 7645 3238
rect 7337 3227 7645 3236
rect 7760 3210 7788 6938
rect 7852 6322 7880 7210
rect 7944 6458 7972 7500
rect 8036 7478 8064 7686
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 8128 6934 8156 8026
rect 8116 6928 8168 6934
rect 8116 6870 8168 6876
rect 8128 6798 8156 6870
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8024 6656 8076 6662
rect 8220 6644 8248 8502
rect 8312 7478 8340 8774
rect 8404 8090 8432 8910
rect 8772 8090 8800 9030
rect 9048 8786 9076 9551
rect 9128 9522 9180 9528
rect 9140 9110 9168 9522
rect 9324 9382 9352 9998
rect 9968 9450 9996 9998
rect 10324 9988 10376 9994
rect 12084 9982 12296 9998
rect 10324 9930 10376 9936
rect 10336 9586 10364 9930
rect 11520 9920 11572 9926
rect 11520 9862 11572 9868
rect 11155 9820 11463 9829
rect 11155 9818 11161 9820
rect 11217 9818 11241 9820
rect 11297 9818 11321 9820
rect 11377 9818 11401 9820
rect 11457 9818 11463 9820
rect 11217 9766 11219 9818
rect 11399 9766 11401 9818
rect 11155 9764 11161 9766
rect 11217 9764 11241 9766
rect 11297 9764 11321 9766
rect 11377 9764 11401 9766
rect 11457 9764 11463 9766
rect 11155 9755 11463 9764
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 9956 9444 10008 9450
rect 9956 9386 10008 9392
rect 10336 9382 10364 9522
rect 11532 9518 11560 9862
rect 10508 9512 10560 9518
rect 10428 9460 10508 9466
rect 10428 9454 10560 9460
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 10428 9438 10548 9454
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 9128 9104 9180 9110
rect 9128 9046 9180 9052
rect 9048 8758 9168 8786
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 8944 8424 8996 8430
rect 8944 8366 8996 8372
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8576 7744 8628 7750
rect 8576 7686 8628 7692
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8300 7472 8352 7478
rect 8300 7414 8352 7420
rect 8024 6598 8076 6604
rect 8128 6616 8248 6644
rect 8300 6656 8352 6662
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 7840 6316 7892 6322
rect 7840 6258 7892 6264
rect 7944 6202 7972 6394
rect 8036 6322 8064 6598
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 7852 6174 7972 6202
rect 7852 5302 7880 6174
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 7944 5710 7972 5850
rect 8036 5846 8064 6258
rect 8024 5840 8076 5846
rect 8024 5782 8076 5788
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 7944 5302 7972 5646
rect 7840 5296 7892 5302
rect 7840 5238 7892 5244
rect 7932 5296 7984 5302
rect 7932 5238 7984 5244
rect 7852 3738 7880 5238
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 7668 3182 7788 3210
rect 7668 3126 7696 3182
rect 7656 3120 7708 3126
rect 7656 3062 7708 3068
rect 7196 2984 7248 2990
rect 7196 2926 7248 2932
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7196 2848 7248 2854
rect 7196 2790 7248 2796
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 7208 2582 7236 2790
rect 7760 2650 7788 2926
rect 7852 2802 7880 3674
rect 7932 2848 7984 2854
rect 7852 2796 7932 2802
rect 7852 2790 7984 2796
rect 7852 2774 7972 2790
rect 8036 2650 8064 5782
rect 8128 3942 8156 6616
rect 8300 6598 8352 6604
rect 8312 6458 8340 6598
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8312 5914 8340 6394
rect 8404 5930 8432 7686
rect 8484 7472 8536 7478
rect 8484 7414 8536 7420
rect 8496 6118 8524 7414
rect 8588 6798 8616 7686
rect 8680 7206 8708 7686
rect 8772 7546 8800 8026
rect 8956 8022 8984 8366
rect 8944 8016 8996 8022
rect 8944 7958 8996 7964
rect 8956 7886 8984 7958
rect 9048 7954 9076 8570
rect 9036 7948 9088 7954
rect 9036 7890 9088 7896
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 9140 7818 9168 8758
rect 9324 8650 9352 9318
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9232 8622 9352 8650
rect 9232 8430 9260 8622
rect 9312 8560 9364 8566
rect 9312 8502 9364 8508
rect 9220 8424 9272 8430
rect 9220 8366 9272 8372
rect 9324 7954 9352 8502
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9588 8016 9640 8022
rect 9588 7958 9640 7964
rect 9312 7948 9364 7954
rect 9312 7890 9364 7896
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 8760 7540 8812 7546
rect 8760 7482 8812 7488
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 8668 7200 8720 7206
rect 8720 7160 8892 7188
rect 8668 7142 8720 7148
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8760 6724 8812 6730
rect 8760 6666 8812 6672
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 8300 5908 8352 5914
rect 8404 5902 8524 5930
rect 8300 5850 8352 5856
rect 8392 5772 8444 5778
rect 8392 5714 8444 5720
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8220 3534 8248 5510
rect 8312 5234 8340 5510
rect 8404 5370 8432 5714
rect 8496 5710 8524 5902
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 8496 5370 8524 5646
rect 8588 5574 8616 5850
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8392 5364 8444 5370
rect 8392 5306 8444 5312
rect 8484 5364 8536 5370
rect 8484 5306 8536 5312
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 8392 5160 8444 5166
rect 8496 5148 8524 5306
rect 8680 5234 8708 6190
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 8444 5120 8524 5148
rect 8392 5102 8444 5108
rect 8772 5030 8800 6666
rect 8864 6390 8892 7160
rect 9048 6458 9076 7482
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9324 6730 9352 7346
rect 9508 6798 9536 7414
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9312 6724 9364 6730
rect 9312 6666 9364 6672
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 8852 6384 8904 6390
rect 8852 6326 8904 6332
rect 9048 5914 9076 6394
rect 9404 6316 9456 6322
rect 9404 6258 9456 6264
rect 9416 6118 9444 6258
rect 9600 6254 9628 7958
rect 9692 7954 9720 8366
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9692 7206 9720 7890
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9692 6934 9720 7142
rect 9680 6928 9732 6934
rect 9680 6870 9732 6876
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9416 5914 9444 6054
rect 9036 5908 9088 5914
rect 9036 5850 9088 5856
rect 9404 5908 9456 5914
rect 9404 5850 9456 5856
rect 9416 5098 9444 5850
rect 9600 5710 9628 6190
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9692 5370 9720 5510
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9404 5092 9456 5098
rect 9404 5034 9456 5040
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 8956 4146 8984 4966
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8300 4004 8352 4010
rect 8300 3946 8352 3952
rect 8312 3738 8340 3946
rect 8956 3942 8984 4082
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9140 3738 9168 3878
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8220 3126 8248 3470
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8208 3120 8260 3126
rect 8484 3120 8536 3126
rect 8208 3062 8260 3068
rect 8404 3080 8484 3108
rect 8404 2922 8432 3080
rect 8484 3062 8536 3068
rect 8588 3058 8616 3130
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 9140 2990 9168 3674
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9324 3126 9352 3334
rect 9312 3120 9364 3126
rect 9312 3062 9364 3068
rect 9128 2984 9180 2990
rect 9128 2926 9180 2932
rect 8392 2916 8444 2922
rect 8392 2858 8444 2864
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 7748 2644 7800 2650
rect 7748 2586 7800 2592
rect 8024 2644 8076 2650
rect 8024 2586 8076 2592
rect 7196 2576 7248 2582
rect 7196 2518 7248 2524
rect 8496 2514 8524 2790
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 8588 2446 8616 2790
rect 9416 2650 9444 5034
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9692 3738 9720 3878
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9784 3058 9812 9114
rect 10428 8634 10456 9438
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 10495 9276 10803 9285
rect 10495 9274 10501 9276
rect 10557 9274 10581 9276
rect 10637 9274 10661 9276
rect 10717 9274 10741 9276
rect 10797 9274 10803 9276
rect 10557 9222 10559 9274
rect 10739 9222 10741 9274
rect 10495 9220 10501 9222
rect 10557 9220 10581 9222
rect 10637 9220 10661 9222
rect 10717 9220 10741 9222
rect 10797 9220 10803 9222
rect 10495 9211 10803 9220
rect 11900 9178 11928 9318
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 12176 9110 12204 9982
rect 12268 9926 12296 9982
rect 12256 9920 12308 9926
rect 12256 9862 12308 9868
rect 13372 9722 13400 10542
rect 13360 9716 13412 9722
rect 13360 9658 13412 9664
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 13188 9178 13216 9522
rect 12256 9172 12308 9178
rect 12256 9114 12308 9120
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 12164 9104 12216 9110
rect 12164 9046 12216 9052
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11155 8732 11463 8741
rect 11155 8730 11161 8732
rect 11217 8730 11241 8732
rect 11297 8730 11321 8732
rect 11377 8730 11401 8732
rect 11457 8730 11463 8732
rect 11217 8678 11219 8730
rect 11399 8678 11401 8730
rect 11155 8676 11161 8678
rect 11217 8676 11241 8678
rect 11297 8676 11321 8678
rect 11377 8676 11401 8678
rect 11457 8676 11463 8678
rect 11155 8667 11463 8676
rect 11532 8634 11560 8910
rect 12164 8900 12216 8906
rect 12164 8842 12216 8848
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11716 8498 11744 8774
rect 12176 8634 12204 8842
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 10060 7546 10088 8434
rect 10495 8188 10803 8197
rect 10495 8186 10501 8188
rect 10557 8186 10581 8188
rect 10637 8186 10661 8188
rect 10717 8186 10741 8188
rect 10797 8186 10803 8188
rect 10557 8134 10559 8186
rect 10739 8134 10741 8186
rect 10495 8132 10501 8134
rect 10557 8132 10581 8134
rect 10637 8132 10661 8134
rect 10717 8132 10741 8134
rect 10797 8132 10803 8134
rect 10495 8123 10803 8132
rect 12268 8090 12296 9114
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12452 7886 12480 8230
rect 13176 7948 13228 7954
rect 13176 7890 13228 7896
rect 12072 7880 12124 7886
rect 12072 7822 12124 7828
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 11155 7644 11463 7653
rect 11155 7642 11161 7644
rect 11217 7642 11241 7644
rect 11297 7642 11321 7644
rect 11377 7642 11401 7644
rect 11457 7642 11463 7644
rect 11217 7590 11219 7642
rect 11399 7590 11401 7642
rect 11155 7588 11161 7590
rect 11217 7588 11241 7590
rect 11297 7588 11321 7590
rect 11377 7588 11401 7590
rect 11457 7588 11463 7590
rect 11155 7579 11463 7588
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 10876 7472 10928 7478
rect 10876 7414 10928 7420
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 10152 7002 10180 7346
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10140 6996 10192 7002
rect 10140 6938 10192 6944
rect 10428 6798 10456 7142
rect 10495 7100 10803 7109
rect 10495 7098 10501 7100
rect 10557 7098 10581 7100
rect 10637 7098 10661 7100
rect 10717 7098 10741 7100
rect 10797 7098 10803 7100
rect 10557 7046 10559 7098
rect 10739 7046 10741 7098
rect 10495 7044 10501 7046
rect 10557 7044 10581 7046
rect 10637 7044 10661 7046
rect 10717 7044 10741 7046
rect 10797 7044 10803 7046
rect 10495 7035 10803 7044
rect 10888 6798 10916 7414
rect 12084 7206 12112 7822
rect 12164 7744 12216 7750
rect 12164 7686 12216 7692
rect 12176 7478 12204 7686
rect 12452 7546 12480 7822
rect 12912 7546 12940 7822
rect 13188 7546 13216 7890
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 12164 7472 12216 7478
rect 12164 7414 12216 7420
rect 13372 7274 13400 7822
rect 13648 7546 13676 9522
rect 13832 7886 13860 11222
rect 14108 11150 14136 11698
rect 14188 11552 14240 11558
rect 14188 11494 14240 11500
rect 14200 11218 14228 11494
rect 14313 11452 14621 11461
rect 14313 11450 14319 11452
rect 14375 11450 14399 11452
rect 14455 11450 14479 11452
rect 14535 11450 14559 11452
rect 14615 11450 14621 11452
rect 14375 11398 14377 11450
rect 14557 11398 14559 11450
rect 14313 11396 14319 11398
rect 14375 11396 14399 11398
rect 14455 11396 14479 11398
rect 14535 11396 14559 11398
rect 14615 11396 14621 11398
rect 14313 11387 14621 11396
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 14844 11150 14872 11698
rect 15028 11354 15056 11698
rect 15200 11688 15252 11694
rect 15200 11630 15252 11636
rect 15212 11354 15240 11630
rect 15016 11348 15068 11354
rect 15016 11290 15068 11296
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 14096 11144 14148 11150
rect 14096 11086 14148 11092
rect 14832 11144 14884 11150
rect 14832 11086 14884 11092
rect 14004 11076 14056 11082
rect 14004 11018 14056 11024
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 12808 7268 12860 7274
rect 12808 7210 12860 7216
rect 13360 7268 13412 7274
rect 13360 7210 13412 7216
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 12084 7002 12112 7142
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10876 6792 10928 6798
rect 10876 6734 10928 6740
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11155 6556 11463 6565
rect 11155 6554 11161 6556
rect 11217 6554 11241 6556
rect 11297 6554 11321 6556
rect 11377 6554 11401 6556
rect 11457 6554 11463 6556
rect 11217 6502 11219 6554
rect 11399 6502 11401 6554
rect 11155 6500 11161 6502
rect 11217 6500 11241 6502
rect 11297 6500 11321 6502
rect 11377 6500 11401 6502
rect 11457 6500 11463 6502
rect 11155 6491 11463 6500
rect 10048 6384 10100 6390
rect 10048 6326 10100 6332
rect 10060 6118 10088 6326
rect 11624 6254 11652 6598
rect 12268 6322 12296 6734
rect 12820 6458 12848 7210
rect 12808 6452 12860 6458
rect 12808 6394 12860 6400
rect 13924 6322 13952 9658
rect 14016 9586 14044 11018
rect 14313 10364 14621 10373
rect 14313 10362 14319 10364
rect 14375 10362 14399 10364
rect 14455 10362 14479 10364
rect 14535 10362 14559 10364
rect 14615 10362 14621 10364
rect 14375 10310 14377 10362
rect 14557 10310 14559 10362
rect 14313 10308 14319 10310
rect 14375 10308 14399 10310
rect 14455 10308 14479 10310
rect 14535 10308 14559 10310
rect 14615 10308 14621 10310
rect 14313 10299 14621 10308
rect 14844 10266 14872 11086
rect 14973 10908 15281 10917
rect 14973 10906 14979 10908
rect 15035 10906 15059 10908
rect 15115 10906 15139 10908
rect 15195 10906 15219 10908
rect 15275 10906 15281 10908
rect 15035 10854 15037 10906
rect 15217 10854 15219 10906
rect 14973 10852 14979 10854
rect 15035 10852 15059 10854
rect 15115 10852 15139 10854
rect 15195 10852 15219 10854
rect 15275 10852 15281 10854
rect 14973 10843 15281 10852
rect 15672 10742 15700 11154
rect 16026 10976 16082 10985
rect 16026 10911 16082 10920
rect 16040 10810 16068 10911
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 15660 10736 15712 10742
rect 15660 10678 15712 10684
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 14832 10056 14884 10062
rect 14832 9998 14884 10004
rect 14004 9580 14056 9586
rect 14004 9522 14056 9528
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 14313 9276 14621 9285
rect 14313 9274 14319 9276
rect 14375 9274 14399 9276
rect 14455 9274 14479 9276
rect 14535 9274 14559 9276
rect 14615 9274 14621 9276
rect 14375 9222 14377 9274
rect 14557 9222 14559 9274
rect 14313 9220 14319 9222
rect 14375 9220 14399 9222
rect 14455 9220 14479 9222
rect 14535 9220 14559 9222
rect 14615 9220 14621 9222
rect 14313 9211 14621 9220
rect 14660 8974 14688 9522
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14752 9178 14780 9454
rect 14844 9178 14872 9998
rect 15660 9988 15712 9994
rect 15660 9930 15712 9936
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 14973 9820 15281 9829
rect 14973 9818 14979 9820
rect 15035 9818 15059 9820
rect 15115 9818 15139 9820
rect 15195 9818 15219 9820
rect 15275 9818 15281 9820
rect 15035 9766 15037 9818
rect 15217 9766 15219 9818
rect 14973 9764 14979 9766
rect 15035 9764 15059 9766
rect 15115 9764 15139 9766
rect 15195 9764 15219 9766
rect 15275 9764 15281 9766
rect 14973 9755 15281 9764
rect 15396 9586 15424 9862
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 14740 9172 14792 9178
rect 14740 9114 14792 9120
rect 14832 9172 14884 9178
rect 14832 9114 14884 9120
rect 14648 8968 14700 8974
rect 14648 8910 14700 8916
rect 14973 8732 15281 8741
rect 14973 8730 14979 8732
rect 15035 8730 15059 8732
rect 15115 8730 15139 8732
rect 15195 8730 15219 8732
rect 15275 8730 15281 8732
rect 15035 8678 15037 8730
rect 15217 8678 15219 8730
rect 14973 8676 14979 8678
rect 15035 8676 15059 8678
rect 15115 8676 15139 8678
rect 15195 8676 15219 8678
rect 15275 8676 15281 8678
rect 14973 8667 15281 8676
rect 15396 8634 15424 9522
rect 15580 9518 15608 9862
rect 15672 9518 15700 9930
rect 16028 9920 16080 9926
rect 16028 9862 16080 9868
rect 16040 9625 16068 9862
rect 16026 9616 16082 9625
rect 16026 9551 16082 9560
rect 15568 9512 15620 9518
rect 15568 9454 15620 9460
rect 15660 9512 15712 9518
rect 15660 9454 15712 9460
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 14313 8188 14621 8197
rect 14313 8186 14319 8188
rect 14375 8186 14399 8188
rect 14455 8186 14479 8188
rect 14535 8186 14559 8188
rect 14615 8186 14621 8188
rect 14375 8134 14377 8186
rect 14557 8134 14559 8186
rect 14313 8132 14319 8134
rect 14375 8132 14399 8134
rect 14455 8132 14479 8134
rect 14535 8132 14559 8134
rect 14615 8132 14621 8134
rect 14313 8123 14621 8132
rect 14372 7948 14424 7954
rect 14372 7890 14424 7896
rect 14384 7546 14412 7890
rect 14752 7886 14780 8434
rect 14832 8424 14884 8430
rect 14832 8366 14884 8372
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14372 7540 14424 7546
rect 14372 7482 14424 7488
rect 14476 7478 14504 7822
rect 14464 7472 14516 7478
rect 14464 7414 14516 7420
rect 14313 7100 14621 7109
rect 14313 7098 14319 7100
rect 14375 7098 14399 7100
rect 14455 7098 14479 7100
rect 14535 7098 14559 7100
rect 14615 7098 14621 7100
rect 14375 7046 14377 7098
rect 14557 7046 14559 7098
rect 14313 7044 14319 7046
rect 14375 7044 14399 7046
rect 14455 7044 14479 7046
rect 14535 7044 14559 7046
rect 14615 7044 14621 7046
rect 14313 7035 14621 7044
rect 14752 6458 14780 7822
rect 14844 7546 14872 8366
rect 14936 8090 14964 8434
rect 14924 8084 14976 8090
rect 14924 8026 14976 8032
rect 15936 7744 15988 7750
rect 15936 7686 15988 7692
rect 14973 7644 15281 7653
rect 14973 7642 14979 7644
rect 15035 7642 15059 7644
rect 15115 7642 15139 7644
rect 15195 7642 15219 7644
rect 15275 7642 15281 7644
rect 15035 7590 15037 7642
rect 15217 7590 15219 7642
rect 14973 7588 14979 7590
rect 15035 7588 15059 7590
rect 15115 7588 15139 7590
rect 15195 7588 15219 7590
rect 15275 7588 15281 7590
rect 14973 7579 15281 7588
rect 15948 7585 15976 7686
rect 15934 7576 15990 7585
rect 14832 7540 14884 7546
rect 15934 7511 15990 7520
rect 14832 7482 14884 7488
rect 14973 6556 15281 6565
rect 14973 6554 14979 6556
rect 15035 6554 15059 6556
rect 15115 6554 15139 6556
rect 15195 6554 15219 6556
rect 15275 6554 15281 6556
rect 15035 6502 15037 6554
rect 15217 6502 15219 6554
rect 14973 6500 14979 6502
rect 15035 6500 15059 6502
rect 15115 6500 15139 6502
rect 15195 6500 15219 6502
rect 15275 6500 15281 6502
rect 14973 6491 15281 6500
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 12256 6316 12308 6322
rect 12256 6258 12308 6264
rect 12900 6316 12952 6322
rect 12900 6258 12952 6264
rect 13912 6316 13964 6322
rect 13912 6258 13964 6264
rect 14556 6316 14608 6322
rect 14740 6316 14792 6322
rect 14608 6276 14688 6304
rect 14556 6258 14608 6264
rect 11612 6248 11664 6254
rect 11612 6190 11664 6196
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 10060 5030 10088 6054
rect 10495 6012 10803 6021
rect 10495 6010 10501 6012
rect 10557 6010 10581 6012
rect 10637 6010 10661 6012
rect 10717 6010 10741 6012
rect 10797 6010 10803 6012
rect 10557 5958 10559 6010
rect 10739 5958 10741 6010
rect 10495 5956 10501 5958
rect 10557 5956 10581 5958
rect 10637 5956 10661 5958
rect 10717 5956 10741 5958
rect 10797 5956 10803 5958
rect 10495 5947 10803 5956
rect 11624 5846 11652 6054
rect 11716 5914 11744 6258
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 11796 6180 11848 6186
rect 11796 6122 11848 6128
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11520 5840 11572 5846
rect 11520 5782 11572 5788
rect 11612 5840 11664 5846
rect 11612 5782 11664 5788
rect 11155 5468 11463 5477
rect 11155 5466 11161 5468
rect 11217 5466 11241 5468
rect 11297 5466 11321 5468
rect 11377 5466 11401 5468
rect 11457 5466 11463 5468
rect 11217 5414 11219 5466
rect 11399 5414 11401 5466
rect 11155 5412 11161 5414
rect 11217 5412 11241 5414
rect 11297 5412 11321 5414
rect 11377 5412 11401 5414
rect 11457 5412 11463 5414
rect 11155 5403 11463 5412
rect 11532 5302 11560 5782
rect 11612 5568 11664 5574
rect 11612 5510 11664 5516
rect 11520 5296 11572 5302
rect 11520 5238 11572 5244
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 10876 5024 10928 5030
rect 10876 4966 10928 4972
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 10428 4826 10456 4966
rect 10495 4924 10803 4933
rect 10495 4922 10501 4924
rect 10557 4922 10581 4924
rect 10637 4922 10661 4924
rect 10717 4922 10741 4924
rect 10797 4922 10803 4924
rect 10557 4870 10559 4922
rect 10739 4870 10741 4922
rect 10495 4868 10501 4870
rect 10557 4868 10581 4870
rect 10637 4868 10661 4870
rect 10717 4868 10741 4870
rect 10797 4868 10803 4870
rect 10495 4859 10803 4868
rect 10888 4826 10916 4966
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 11256 4758 11284 4966
rect 11624 4826 11652 5510
rect 11716 5302 11744 5850
rect 11808 5710 11836 6122
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 11992 5914 12020 6054
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 12452 5574 12480 6190
rect 12912 5710 12940 6258
rect 12992 6248 13044 6254
rect 12992 6190 13044 6196
rect 13004 5914 13032 6190
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 12900 5704 12952 5710
rect 12900 5646 12952 5652
rect 12440 5568 12492 5574
rect 12440 5510 12492 5516
rect 11704 5296 11756 5302
rect 11704 5238 11756 5244
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11612 4820 11664 4826
rect 11612 4762 11664 4768
rect 11244 4752 11296 4758
rect 11244 4694 11296 4700
rect 11060 4684 11112 4690
rect 11060 4626 11112 4632
rect 11072 4146 11100 4626
rect 11155 4380 11463 4389
rect 11155 4378 11161 4380
rect 11217 4378 11241 4380
rect 11297 4378 11321 4380
rect 11377 4378 11401 4380
rect 11457 4378 11463 4380
rect 11217 4326 11219 4378
rect 11399 4326 11401 4378
rect 11155 4324 11161 4326
rect 11217 4324 11241 4326
rect 11297 4324 11321 4326
rect 11377 4324 11401 4326
rect 11457 4324 11463 4326
rect 11155 4315 11463 4324
rect 11900 4146 11928 4966
rect 12912 4146 12940 5646
rect 13004 5234 13032 5850
rect 13924 5710 13952 6258
rect 14096 6112 14148 6118
rect 14096 6054 14148 6060
rect 14108 5778 14136 6054
rect 14313 6012 14621 6021
rect 14313 6010 14319 6012
rect 14375 6010 14399 6012
rect 14455 6010 14479 6012
rect 14535 6010 14559 6012
rect 14615 6010 14621 6012
rect 14375 5958 14377 6010
rect 14557 5958 14559 6010
rect 14313 5956 14319 5958
rect 14375 5956 14399 5958
rect 14455 5956 14479 5958
rect 14535 5956 14559 5958
rect 14615 5956 14621 5958
rect 14313 5947 14621 5956
rect 14660 5914 14688 6276
rect 14740 6258 14792 6264
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 14096 5772 14148 5778
rect 14096 5714 14148 5720
rect 14752 5710 14780 6258
rect 13360 5704 13412 5710
rect 13360 5646 13412 5652
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 13176 5568 13228 5574
rect 13176 5510 13228 5516
rect 13188 5234 13216 5510
rect 13372 5370 13400 5646
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 14313 4924 14621 4933
rect 14313 4922 14319 4924
rect 14375 4922 14399 4924
rect 14455 4922 14479 4924
rect 14535 4922 14559 4924
rect 14615 4922 14621 4924
rect 14375 4870 14377 4922
rect 14557 4870 14559 4922
rect 14313 4868 14319 4870
rect 14375 4868 14399 4870
rect 14455 4868 14479 4870
rect 14535 4868 14559 4870
rect 14615 4868 14621 4870
rect 14313 4859 14621 4868
rect 14752 4146 14780 5646
rect 16028 5568 16080 5574
rect 16026 5536 16028 5545
rect 16080 5536 16082 5545
rect 14973 5468 15281 5477
rect 16026 5471 16082 5480
rect 14973 5466 14979 5468
rect 15035 5466 15059 5468
rect 15115 5466 15139 5468
rect 15195 5466 15219 5468
rect 15275 5466 15281 5468
rect 15035 5414 15037 5466
rect 15217 5414 15219 5466
rect 14973 5412 14979 5414
rect 15035 5412 15059 5414
rect 15115 5412 15139 5414
rect 15195 5412 15219 5414
rect 15275 5412 15281 5414
rect 14973 5403 15281 5412
rect 14973 4380 15281 4389
rect 14973 4378 14979 4380
rect 15035 4378 15059 4380
rect 15115 4378 15139 4380
rect 15195 4378 15219 4380
rect 15275 4378 15281 4380
rect 15035 4326 15037 4378
rect 15217 4326 15219 4378
rect 14973 4324 14979 4326
rect 15035 4324 15059 4326
rect 15115 4324 15139 4326
rect 15195 4324 15219 4326
rect 15275 4324 15281 4326
rect 14973 4315 15281 4324
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 12532 4004 12584 4010
rect 12532 3946 12584 3952
rect 10495 3836 10803 3845
rect 10495 3834 10501 3836
rect 10557 3834 10581 3836
rect 10637 3834 10661 3836
rect 10717 3834 10741 3836
rect 10797 3834 10803 3836
rect 10557 3782 10559 3834
rect 10739 3782 10741 3834
rect 10495 3780 10501 3782
rect 10557 3780 10581 3782
rect 10637 3780 10661 3782
rect 10717 3780 10741 3782
rect 10797 3780 10803 3782
rect 10495 3771 10803 3780
rect 12544 3534 12572 3946
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 12636 3602 12664 3878
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 13556 3534 13584 3878
rect 13740 3738 13768 4082
rect 14016 3738 14044 4082
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 14108 3466 14136 4082
rect 14313 3836 14621 3845
rect 14313 3834 14319 3836
rect 14375 3834 14399 3836
rect 14455 3834 14479 3836
rect 14535 3834 14559 3836
rect 14615 3834 14621 3836
rect 14375 3782 14377 3834
rect 14557 3782 14559 3834
rect 14313 3780 14319 3782
rect 14375 3780 14399 3782
rect 14455 3780 14479 3782
rect 14535 3780 14559 3782
rect 14615 3780 14621 3782
rect 14313 3771 14621 3780
rect 15936 3664 15988 3670
rect 15936 3606 15988 3612
rect 15948 3505 15976 3606
rect 15934 3496 15990 3505
rect 14096 3460 14148 3466
rect 15934 3431 15990 3440
rect 14096 3402 14148 3408
rect 13176 3392 13228 3398
rect 13176 3334 13228 3340
rect 11155 3292 11463 3301
rect 11155 3290 11161 3292
rect 11217 3290 11241 3292
rect 11297 3290 11321 3292
rect 11377 3290 11401 3292
rect 11457 3290 11463 3292
rect 11217 3238 11219 3290
rect 11399 3238 11401 3290
rect 11155 3236 11161 3238
rect 11217 3236 11241 3238
rect 11297 3236 11321 3238
rect 11377 3236 11401 3238
rect 11457 3236 11463 3238
rect 11155 3227 11463 3236
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 9784 2774 9812 2994
rect 10416 2984 10468 2990
rect 10416 2926 10468 2932
rect 11428 2984 11480 2990
rect 11612 2984 11664 2990
rect 11480 2944 11612 2972
rect 11428 2926 11480 2932
rect 11612 2926 11664 2932
rect 9784 2746 9996 2774
rect 9404 2644 9456 2650
rect 9404 2586 9456 2592
rect 9968 2446 9996 2746
rect 10428 2446 10456 2926
rect 12440 2916 12492 2922
rect 12440 2858 12492 2864
rect 10876 2848 10928 2854
rect 10876 2790 10928 2796
rect 10495 2748 10803 2757
rect 10495 2746 10501 2748
rect 10557 2746 10581 2748
rect 10637 2746 10661 2748
rect 10717 2746 10741 2748
rect 10797 2746 10803 2748
rect 10557 2694 10559 2746
rect 10739 2694 10741 2746
rect 10495 2692 10501 2694
rect 10557 2692 10581 2694
rect 10637 2692 10661 2694
rect 10717 2692 10741 2694
rect 10797 2692 10803 2694
rect 10495 2683 10803 2692
rect 10888 2650 10916 2790
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 12452 2446 12480 2858
rect 13188 2854 13216 3334
rect 14973 3292 15281 3301
rect 14973 3290 14979 3292
rect 15035 3290 15059 3292
rect 15115 3290 15139 3292
rect 15195 3290 15219 3292
rect 15275 3290 15281 3292
rect 15035 3238 15037 3290
rect 15217 3238 15219 3290
rect 14973 3236 14979 3238
rect 15035 3236 15059 3238
rect 15115 3236 15139 3238
rect 15195 3236 15219 3238
rect 15275 3236 15281 3238
rect 14973 3227 15281 3236
rect 13176 2848 13228 2854
rect 13176 2790 13228 2796
rect 14313 2748 14621 2757
rect 14313 2746 14319 2748
rect 14375 2746 14399 2748
rect 14455 2746 14479 2748
rect 14535 2746 14559 2748
rect 14615 2746 14621 2748
rect 14375 2694 14377 2746
rect 14557 2694 14559 2746
rect 14313 2692 14319 2694
rect 14375 2692 14399 2694
rect 14455 2692 14479 2694
rect 14535 2692 14559 2694
rect 14615 2692 14621 2694
rect 14313 2683 14621 2692
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 10416 2440 10468 2446
rect 12440 2440 12492 2446
rect 10416 2382 10468 2388
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 3519 2204 3827 2213
rect 3519 2202 3525 2204
rect 3581 2202 3605 2204
rect 3661 2202 3685 2204
rect 3741 2202 3765 2204
rect 3821 2202 3827 2204
rect 3581 2150 3583 2202
rect 3763 2150 3765 2202
rect 3519 2148 3525 2150
rect 3581 2148 3605 2150
rect 3661 2148 3685 2150
rect 3741 2148 3765 2150
rect 3821 2148 3827 2150
rect 3519 2139 3827 2148
rect 4540 800 4568 2246
rect 7208 1306 7236 2382
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 7337 2204 7645 2213
rect 7337 2202 7343 2204
rect 7399 2202 7423 2204
rect 7479 2202 7503 2204
rect 7559 2202 7583 2204
rect 7639 2202 7645 2204
rect 7399 2150 7401 2202
rect 7581 2150 7583 2202
rect 7337 2148 7343 2150
rect 7399 2148 7423 2150
rect 7479 2148 7503 2150
rect 7559 2148 7583 2150
rect 7639 2148 7645 2150
rect 7337 2139 7645 2148
rect 7116 1278 7236 1306
rect 7116 800 7144 1278
rect 7760 800 7788 2246
rect 8404 800 8432 2246
rect 9140 1306 9168 2382
rect 12268 2366 12388 2394
rect 12440 2382 12492 2388
rect 11155 2204 11463 2213
rect 11155 2202 11161 2204
rect 11217 2202 11241 2204
rect 11297 2202 11321 2204
rect 11377 2202 11401 2204
rect 11457 2202 11463 2204
rect 11217 2150 11219 2202
rect 11399 2150 11401 2202
rect 11155 2148 11161 2150
rect 11217 2148 11241 2150
rect 11297 2148 11321 2150
rect 11377 2148 11401 2150
rect 11457 2148 11463 2150
rect 11155 2139 11463 2148
rect 9048 1278 9168 1306
rect 9048 800 9076 1278
rect 12268 800 12296 2366
rect 12360 2310 12388 2366
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 14973 2204 15281 2213
rect 14973 2202 14979 2204
rect 15035 2202 15059 2204
rect 15115 2202 15139 2204
rect 15195 2202 15219 2204
rect 15275 2202 15281 2204
rect 15035 2150 15037 2202
rect 15217 2150 15219 2202
rect 14973 2148 14979 2150
rect 15035 2148 15059 2150
rect 15115 2148 15139 2150
rect 15195 2148 15219 2150
rect 15275 2148 15281 2150
rect 14973 2139 15281 2148
rect 4526 0 4582 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 12254 0 12310 800
<< via2 >>
rect 3525 17434 3581 17436
rect 3605 17434 3661 17436
rect 3685 17434 3741 17436
rect 3765 17434 3821 17436
rect 3525 17382 3571 17434
rect 3571 17382 3581 17434
rect 3605 17382 3635 17434
rect 3635 17382 3647 17434
rect 3647 17382 3661 17434
rect 3685 17382 3699 17434
rect 3699 17382 3711 17434
rect 3711 17382 3741 17434
rect 3765 17382 3775 17434
rect 3775 17382 3821 17434
rect 3525 17380 3581 17382
rect 3605 17380 3661 17382
rect 3685 17380 3741 17382
rect 3765 17380 3821 17382
rect 7343 17434 7399 17436
rect 7423 17434 7479 17436
rect 7503 17434 7559 17436
rect 7583 17434 7639 17436
rect 7343 17382 7389 17434
rect 7389 17382 7399 17434
rect 7423 17382 7453 17434
rect 7453 17382 7465 17434
rect 7465 17382 7479 17434
rect 7503 17382 7517 17434
rect 7517 17382 7529 17434
rect 7529 17382 7559 17434
rect 7583 17382 7593 17434
rect 7593 17382 7639 17434
rect 7343 17380 7399 17382
rect 7423 17380 7479 17382
rect 7503 17380 7559 17382
rect 7583 17380 7639 17382
rect 11161 17434 11217 17436
rect 11241 17434 11297 17436
rect 11321 17434 11377 17436
rect 11401 17434 11457 17436
rect 11161 17382 11207 17434
rect 11207 17382 11217 17434
rect 11241 17382 11271 17434
rect 11271 17382 11283 17434
rect 11283 17382 11297 17434
rect 11321 17382 11335 17434
rect 11335 17382 11347 17434
rect 11347 17382 11377 17434
rect 11401 17382 11411 17434
rect 11411 17382 11457 17434
rect 11161 17380 11217 17382
rect 11241 17380 11297 17382
rect 11321 17380 11377 17382
rect 11401 17380 11457 17382
rect 14979 17434 15035 17436
rect 15059 17434 15115 17436
rect 15139 17434 15195 17436
rect 15219 17434 15275 17436
rect 14979 17382 15025 17434
rect 15025 17382 15035 17434
rect 15059 17382 15089 17434
rect 15089 17382 15101 17434
rect 15101 17382 15115 17434
rect 15139 17382 15153 17434
rect 15153 17382 15165 17434
rect 15165 17382 15195 17434
rect 15219 17382 15229 17434
rect 15229 17382 15275 17434
rect 14979 17380 15035 17382
rect 15059 17380 15115 17382
rect 15139 17380 15195 17382
rect 15219 17380 15275 17382
rect 2865 16890 2921 16892
rect 2945 16890 3001 16892
rect 3025 16890 3081 16892
rect 3105 16890 3161 16892
rect 2865 16838 2911 16890
rect 2911 16838 2921 16890
rect 2945 16838 2975 16890
rect 2975 16838 2987 16890
rect 2987 16838 3001 16890
rect 3025 16838 3039 16890
rect 3039 16838 3051 16890
rect 3051 16838 3081 16890
rect 3105 16838 3115 16890
rect 3115 16838 3161 16890
rect 2865 16836 2921 16838
rect 2945 16836 3001 16838
rect 3025 16836 3081 16838
rect 3105 16836 3161 16838
rect 6683 16890 6739 16892
rect 6763 16890 6819 16892
rect 6843 16890 6899 16892
rect 6923 16890 6979 16892
rect 6683 16838 6729 16890
rect 6729 16838 6739 16890
rect 6763 16838 6793 16890
rect 6793 16838 6805 16890
rect 6805 16838 6819 16890
rect 6843 16838 6857 16890
rect 6857 16838 6869 16890
rect 6869 16838 6899 16890
rect 6923 16838 6933 16890
rect 6933 16838 6979 16890
rect 6683 16836 6739 16838
rect 6763 16836 6819 16838
rect 6843 16836 6899 16838
rect 6923 16836 6979 16838
rect 3525 16346 3581 16348
rect 3605 16346 3661 16348
rect 3685 16346 3741 16348
rect 3765 16346 3821 16348
rect 3525 16294 3571 16346
rect 3571 16294 3581 16346
rect 3605 16294 3635 16346
rect 3635 16294 3647 16346
rect 3647 16294 3661 16346
rect 3685 16294 3699 16346
rect 3699 16294 3711 16346
rect 3711 16294 3741 16346
rect 3765 16294 3775 16346
rect 3775 16294 3821 16346
rect 3525 16292 3581 16294
rect 3605 16292 3661 16294
rect 3685 16292 3741 16294
rect 3765 16292 3821 16294
rect 2865 15802 2921 15804
rect 2945 15802 3001 15804
rect 3025 15802 3081 15804
rect 3105 15802 3161 15804
rect 2865 15750 2911 15802
rect 2911 15750 2921 15802
rect 2945 15750 2975 15802
rect 2975 15750 2987 15802
rect 2987 15750 3001 15802
rect 3025 15750 3039 15802
rect 3039 15750 3051 15802
rect 3051 15750 3081 15802
rect 3105 15750 3115 15802
rect 3115 15750 3161 15802
rect 2865 15748 2921 15750
rect 2945 15748 3001 15750
rect 3025 15748 3081 15750
rect 3105 15748 3161 15750
rect 3525 15258 3581 15260
rect 3605 15258 3661 15260
rect 3685 15258 3741 15260
rect 3765 15258 3821 15260
rect 3525 15206 3571 15258
rect 3571 15206 3581 15258
rect 3605 15206 3635 15258
rect 3635 15206 3647 15258
rect 3647 15206 3661 15258
rect 3685 15206 3699 15258
rect 3699 15206 3711 15258
rect 3711 15206 3741 15258
rect 3765 15206 3775 15258
rect 3775 15206 3821 15258
rect 3525 15204 3581 15206
rect 3605 15204 3661 15206
rect 3685 15204 3741 15206
rect 3765 15204 3821 15206
rect 938 14340 994 14376
rect 938 14320 940 14340
rect 940 14320 992 14340
rect 992 14320 994 14340
rect 938 12960 994 13016
rect 1398 12280 1454 12336
rect 1398 10920 1454 10976
rect 938 10240 994 10296
rect 1490 9560 1546 9616
rect 938 8900 994 8936
rect 938 8880 940 8900
rect 940 8880 992 8900
rect 992 8880 994 8900
rect 938 7520 994 7576
rect 2865 14714 2921 14716
rect 2945 14714 3001 14716
rect 3025 14714 3081 14716
rect 3105 14714 3161 14716
rect 2865 14662 2911 14714
rect 2911 14662 2921 14714
rect 2945 14662 2975 14714
rect 2975 14662 2987 14714
rect 2987 14662 3001 14714
rect 3025 14662 3039 14714
rect 3039 14662 3051 14714
rect 3051 14662 3081 14714
rect 3105 14662 3115 14714
rect 3115 14662 3161 14714
rect 2865 14660 2921 14662
rect 2945 14660 3001 14662
rect 3025 14660 3081 14662
rect 3105 14660 3161 14662
rect 6683 15802 6739 15804
rect 6763 15802 6819 15804
rect 6843 15802 6899 15804
rect 6923 15802 6979 15804
rect 6683 15750 6729 15802
rect 6729 15750 6739 15802
rect 6763 15750 6793 15802
rect 6793 15750 6805 15802
rect 6805 15750 6819 15802
rect 6843 15750 6857 15802
rect 6857 15750 6869 15802
rect 6869 15750 6899 15802
rect 6923 15750 6933 15802
rect 6933 15750 6979 15802
rect 6683 15748 6739 15750
rect 6763 15748 6819 15750
rect 6843 15748 6899 15750
rect 6923 15748 6979 15750
rect 7343 16346 7399 16348
rect 7423 16346 7479 16348
rect 7503 16346 7559 16348
rect 7583 16346 7639 16348
rect 7343 16294 7389 16346
rect 7389 16294 7399 16346
rect 7423 16294 7453 16346
rect 7453 16294 7465 16346
rect 7465 16294 7479 16346
rect 7503 16294 7517 16346
rect 7517 16294 7529 16346
rect 7529 16294 7559 16346
rect 7583 16294 7593 16346
rect 7593 16294 7639 16346
rect 7343 16292 7399 16294
rect 7423 16292 7479 16294
rect 7503 16292 7559 16294
rect 7583 16292 7639 16294
rect 3525 14170 3581 14172
rect 3605 14170 3661 14172
rect 3685 14170 3741 14172
rect 3765 14170 3821 14172
rect 3525 14118 3571 14170
rect 3571 14118 3581 14170
rect 3605 14118 3635 14170
rect 3635 14118 3647 14170
rect 3647 14118 3661 14170
rect 3685 14118 3699 14170
rect 3699 14118 3711 14170
rect 3711 14118 3741 14170
rect 3765 14118 3775 14170
rect 3775 14118 3821 14170
rect 3525 14116 3581 14118
rect 3605 14116 3661 14118
rect 3685 14116 3741 14118
rect 3765 14116 3821 14118
rect 2865 13626 2921 13628
rect 2945 13626 3001 13628
rect 3025 13626 3081 13628
rect 3105 13626 3161 13628
rect 2865 13574 2911 13626
rect 2911 13574 2921 13626
rect 2945 13574 2975 13626
rect 2975 13574 2987 13626
rect 2987 13574 3001 13626
rect 3025 13574 3039 13626
rect 3039 13574 3051 13626
rect 3051 13574 3081 13626
rect 3105 13574 3115 13626
rect 3115 13574 3161 13626
rect 2865 13572 2921 13574
rect 2945 13572 3001 13574
rect 3025 13572 3081 13574
rect 3105 13572 3161 13574
rect 3525 13082 3581 13084
rect 3605 13082 3661 13084
rect 3685 13082 3741 13084
rect 3765 13082 3821 13084
rect 3525 13030 3571 13082
rect 3571 13030 3581 13082
rect 3605 13030 3635 13082
rect 3635 13030 3647 13082
rect 3647 13030 3661 13082
rect 3685 13030 3699 13082
rect 3699 13030 3711 13082
rect 3711 13030 3741 13082
rect 3765 13030 3775 13082
rect 3775 13030 3821 13082
rect 3525 13028 3581 13030
rect 3605 13028 3661 13030
rect 3685 13028 3741 13030
rect 3765 13028 3821 13030
rect 2865 12538 2921 12540
rect 2945 12538 3001 12540
rect 3025 12538 3081 12540
rect 3105 12538 3161 12540
rect 2865 12486 2911 12538
rect 2911 12486 2921 12538
rect 2945 12486 2975 12538
rect 2975 12486 2987 12538
rect 2987 12486 3001 12538
rect 3025 12486 3039 12538
rect 3039 12486 3051 12538
rect 3051 12486 3081 12538
rect 3105 12486 3115 12538
rect 3115 12486 3161 12538
rect 2865 12484 2921 12486
rect 2945 12484 3001 12486
rect 3025 12484 3081 12486
rect 3105 12484 3161 12486
rect 3525 11994 3581 11996
rect 3605 11994 3661 11996
rect 3685 11994 3741 11996
rect 3765 11994 3821 11996
rect 3525 11942 3571 11994
rect 3571 11942 3581 11994
rect 3605 11942 3635 11994
rect 3635 11942 3647 11994
rect 3647 11942 3661 11994
rect 3685 11942 3699 11994
rect 3699 11942 3711 11994
rect 3711 11942 3741 11994
rect 3765 11942 3775 11994
rect 3775 11942 3821 11994
rect 3525 11940 3581 11942
rect 3605 11940 3661 11942
rect 3685 11940 3741 11942
rect 3765 11940 3821 11942
rect 2865 11450 2921 11452
rect 2945 11450 3001 11452
rect 3025 11450 3081 11452
rect 3105 11450 3161 11452
rect 2865 11398 2911 11450
rect 2911 11398 2921 11450
rect 2945 11398 2975 11450
rect 2975 11398 2987 11450
rect 2987 11398 3001 11450
rect 3025 11398 3039 11450
rect 3039 11398 3051 11450
rect 3051 11398 3081 11450
rect 3105 11398 3115 11450
rect 3115 11398 3161 11450
rect 2865 11396 2921 11398
rect 2945 11396 3001 11398
rect 3025 11396 3081 11398
rect 3105 11396 3161 11398
rect 3525 10906 3581 10908
rect 3605 10906 3661 10908
rect 3685 10906 3741 10908
rect 3765 10906 3821 10908
rect 3525 10854 3571 10906
rect 3571 10854 3581 10906
rect 3605 10854 3635 10906
rect 3635 10854 3647 10906
rect 3647 10854 3661 10906
rect 3685 10854 3699 10906
rect 3699 10854 3711 10906
rect 3711 10854 3741 10906
rect 3765 10854 3775 10906
rect 3775 10854 3821 10906
rect 3525 10852 3581 10854
rect 3605 10852 3661 10854
rect 3685 10852 3741 10854
rect 3765 10852 3821 10854
rect 2865 10362 2921 10364
rect 2945 10362 3001 10364
rect 3025 10362 3081 10364
rect 3105 10362 3161 10364
rect 2865 10310 2911 10362
rect 2911 10310 2921 10362
rect 2945 10310 2975 10362
rect 2975 10310 2987 10362
rect 2987 10310 3001 10362
rect 3025 10310 3039 10362
rect 3039 10310 3051 10362
rect 3051 10310 3081 10362
rect 3105 10310 3115 10362
rect 3115 10310 3161 10362
rect 2865 10308 2921 10310
rect 2945 10308 3001 10310
rect 3025 10308 3081 10310
rect 3105 10308 3161 10310
rect 3525 9818 3581 9820
rect 3605 9818 3661 9820
rect 3685 9818 3741 9820
rect 3765 9818 3821 9820
rect 3525 9766 3571 9818
rect 3571 9766 3581 9818
rect 3605 9766 3635 9818
rect 3635 9766 3647 9818
rect 3647 9766 3661 9818
rect 3685 9766 3699 9818
rect 3699 9766 3711 9818
rect 3711 9766 3741 9818
rect 3765 9766 3775 9818
rect 3775 9766 3821 9818
rect 3525 9764 3581 9766
rect 3605 9764 3661 9766
rect 3685 9764 3741 9766
rect 3765 9764 3821 9766
rect 2865 9274 2921 9276
rect 2945 9274 3001 9276
rect 3025 9274 3081 9276
rect 3105 9274 3161 9276
rect 2865 9222 2911 9274
rect 2911 9222 2921 9274
rect 2945 9222 2975 9274
rect 2975 9222 2987 9274
rect 2987 9222 3001 9274
rect 3025 9222 3039 9274
rect 3039 9222 3051 9274
rect 3051 9222 3081 9274
rect 3105 9222 3115 9274
rect 3115 9222 3161 9274
rect 2865 9220 2921 9222
rect 2945 9220 3001 9222
rect 3025 9220 3081 9222
rect 3105 9220 3161 9222
rect 3525 8730 3581 8732
rect 3605 8730 3661 8732
rect 3685 8730 3741 8732
rect 3765 8730 3821 8732
rect 3525 8678 3571 8730
rect 3571 8678 3581 8730
rect 3605 8678 3635 8730
rect 3635 8678 3647 8730
rect 3647 8678 3661 8730
rect 3685 8678 3699 8730
rect 3699 8678 3711 8730
rect 3711 8678 3741 8730
rect 3765 8678 3775 8730
rect 3775 8678 3821 8730
rect 3525 8676 3581 8678
rect 3605 8676 3661 8678
rect 3685 8676 3741 8678
rect 3765 8676 3821 8678
rect 2686 8200 2742 8256
rect 2865 8186 2921 8188
rect 2945 8186 3001 8188
rect 3025 8186 3081 8188
rect 3105 8186 3161 8188
rect 2865 8134 2911 8186
rect 2911 8134 2921 8186
rect 2945 8134 2975 8186
rect 2975 8134 2987 8186
rect 2987 8134 3001 8186
rect 3025 8134 3039 8186
rect 3039 8134 3051 8186
rect 3051 8134 3081 8186
rect 3105 8134 3115 8186
rect 3115 8134 3161 8186
rect 2865 8132 2921 8134
rect 2945 8132 3001 8134
rect 3025 8132 3081 8134
rect 3105 8132 3161 8134
rect 2502 7792 2558 7848
rect 938 6840 994 6896
rect 938 5480 994 5536
rect 1398 4664 1454 4720
rect 1030 4156 1032 4176
rect 1032 4156 1084 4176
rect 1084 4156 1086 4176
rect 1030 4120 1086 4156
rect 938 3476 940 3496
rect 940 3476 992 3496
rect 992 3476 994 3496
rect 938 3440 994 3476
rect 2865 7098 2921 7100
rect 2945 7098 3001 7100
rect 3025 7098 3081 7100
rect 3105 7098 3161 7100
rect 2865 7046 2911 7098
rect 2911 7046 2921 7098
rect 2945 7046 2975 7098
rect 2975 7046 2987 7098
rect 2987 7046 3001 7098
rect 3025 7046 3039 7098
rect 3039 7046 3051 7098
rect 3051 7046 3081 7098
rect 3105 7046 3115 7098
rect 3115 7046 3161 7098
rect 2865 7044 2921 7046
rect 2945 7044 3001 7046
rect 3025 7044 3081 7046
rect 3105 7044 3161 7046
rect 2778 6160 2834 6216
rect 2865 6010 2921 6012
rect 2945 6010 3001 6012
rect 3025 6010 3081 6012
rect 3105 6010 3161 6012
rect 2865 5958 2911 6010
rect 2911 5958 2921 6010
rect 2945 5958 2975 6010
rect 2975 5958 2987 6010
rect 2987 5958 3001 6010
rect 3025 5958 3039 6010
rect 3039 5958 3051 6010
rect 3051 5958 3081 6010
rect 3105 5958 3115 6010
rect 3115 5958 3161 6010
rect 2865 5956 2921 5958
rect 2945 5956 3001 5958
rect 3025 5956 3081 5958
rect 3105 5956 3161 5958
rect 3525 7642 3581 7644
rect 3605 7642 3661 7644
rect 3685 7642 3741 7644
rect 3765 7642 3821 7644
rect 3525 7590 3571 7642
rect 3571 7590 3581 7642
rect 3605 7590 3635 7642
rect 3635 7590 3647 7642
rect 3647 7590 3661 7642
rect 3685 7590 3699 7642
rect 3699 7590 3711 7642
rect 3711 7590 3741 7642
rect 3765 7590 3775 7642
rect 3775 7590 3821 7642
rect 3525 7588 3581 7590
rect 3605 7588 3661 7590
rect 3685 7588 3741 7590
rect 3765 7588 3821 7590
rect 7343 15258 7399 15260
rect 7423 15258 7479 15260
rect 7503 15258 7559 15260
rect 7583 15258 7639 15260
rect 7343 15206 7389 15258
rect 7389 15206 7399 15258
rect 7423 15206 7453 15258
rect 7453 15206 7465 15258
rect 7465 15206 7479 15258
rect 7503 15206 7517 15258
rect 7517 15206 7529 15258
rect 7529 15206 7559 15258
rect 7583 15206 7593 15258
rect 7593 15206 7639 15258
rect 7343 15204 7399 15206
rect 7423 15204 7479 15206
rect 7503 15204 7559 15206
rect 7583 15204 7639 15206
rect 6683 14714 6739 14716
rect 6763 14714 6819 14716
rect 6843 14714 6899 14716
rect 6923 14714 6979 14716
rect 6683 14662 6729 14714
rect 6729 14662 6739 14714
rect 6763 14662 6793 14714
rect 6793 14662 6805 14714
rect 6805 14662 6819 14714
rect 6843 14662 6857 14714
rect 6857 14662 6869 14714
rect 6869 14662 6899 14714
rect 6923 14662 6933 14714
rect 6933 14662 6979 14714
rect 6683 14660 6739 14662
rect 6763 14660 6819 14662
rect 6843 14660 6899 14662
rect 6923 14660 6979 14662
rect 6683 13626 6739 13628
rect 6763 13626 6819 13628
rect 6843 13626 6899 13628
rect 6923 13626 6979 13628
rect 6683 13574 6729 13626
rect 6729 13574 6739 13626
rect 6763 13574 6793 13626
rect 6793 13574 6805 13626
rect 6805 13574 6819 13626
rect 6843 13574 6857 13626
rect 6857 13574 6869 13626
rect 6869 13574 6899 13626
rect 6923 13574 6933 13626
rect 6933 13574 6979 13626
rect 6683 13572 6739 13574
rect 6763 13572 6819 13574
rect 6843 13572 6899 13574
rect 6923 13572 6979 13574
rect 7343 14170 7399 14172
rect 7423 14170 7479 14172
rect 7503 14170 7559 14172
rect 7583 14170 7639 14172
rect 7343 14118 7389 14170
rect 7389 14118 7399 14170
rect 7423 14118 7453 14170
rect 7453 14118 7465 14170
rect 7465 14118 7479 14170
rect 7503 14118 7517 14170
rect 7517 14118 7529 14170
rect 7529 14118 7559 14170
rect 7583 14118 7593 14170
rect 7593 14118 7639 14170
rect 7343 14116 7399 14118
rect 7423 14116 7479 14118
rect 7503 14116 7559 14118
rect 7583 14116 7639 14118
rect 4342 7828 4344 7848
rect 4344 7828 4396 7848
rect 4396 7828 4398 7848
rect 4342 7792 4398 7828
rect 4250 7284 4252 7304
rect 4252 7284 4304 7304
rect 4304 7284 4306 7304
rect 4250 7248 4306 7284
rect 3525 6554 3581 6556
rect 3605 6554 3661 6556
rect 3685 6554 3741 6556
rect 3765 6554 3821 6556
rect 3525 6502 3571 6554
rect 3571 6502 3581 6554
rect 3605 6502 3635 6554
rect 3635 6502 3647 6554
rect 3647 6502 3661 6554
rect 3685 6502 3699 6554
rect 3699 6502 3711 6554
rect 3711 6502 3741 6554
rect 3765 6502 3775 6554
rect 3775 6502 3821 6554
rect 3525 6500 3581 6502
rect 3605 6500 3661 6502
rect 3685 6500 3741 6502
rect 3765 6500 3821 6502
rect 2865 4922 2921 4924
rect 2945 4922 3001 4924
rect 3025 4922 3081 4924
rect 3105 4922 3161 4924
rect 2865 4870 2911 4922
rect 2911 4870 2921 4922
rect 2945 4870 2975 4922
rect 2975 4870 2987 4922
rect 2987 4870 3001 4922
rect 3025 4870 3039 4922
rect 3039 4870 3051 4922
rect 3051 4870 3081 4922
rect 3105 4870 3115 4922
rect 3115 4870 3161 4922
rect 2865 4868 2921 4870
rect 2945 4868 3001 4870
rect 3025 4868 3081 4870
rect 3105 4868 3161 4870
rect 2865 3834 2921 3836
rect 2945 3834 3001 3836
rect 3025 3834 3081 3836
rect 3105 3834 3161 3836
rect 2865 3782 2911 3834
rect 2911 3782 2921 3834
rect 2945 3782 2975 3834
rect 2975 3782 2987 3834
rect 2987 3782 3001 3834
rect 3025 3782 3039 3834
rect 3039 3782 3051 3834
rect 3051 3782 3081 3834
rect 3105 3782 3115 3834
rect 3115 3782 3161 3834
rect 2865 3780 2921 3782
rect 2945 3780 3001 3782
rect 3025 3780 3081 3782
rect 3105 3780 3161 3782
rect 3525 5466 3581 5468
rect 3605 5466 3661 5468
rect 3685 5466 3741 5468
rect 3765 5466 3821 5468
rect 3525 5414 3571 5466
rect 3571 5414 3581 5466
rect 3605 5414 3635 5466
rect 3635 5414 3647 5466
rect 3647 5414 3661 5466
rect 3685 5414 3699 5466
rect 3699 5414 3711 5466
rect 3711 5414 3741 5466
rect 3765 5414 3775 5466
rect 3775 5414 3821 5466
rect 3525 5412 3581 5414
rect 3605 5412 3661 5414
rect 3685 5412 3741 5414
rect 3765 5412 3821 5414
rect 3525 4378 3581 4380
rect 3605 4378 3661 4380
rect 3685 4378 3741 4380
rect 3765 4378 3821 4380
rect 3525 4326 3571 4378
rect 3571 4326 3581 4378
rect 3605 4326 3635 4378
rect 3635 4326 3647 4378
rect 3647 4326 3661 4378
rect 3685 4326 3699 4378
rect 3699 4326 3711 4378
rect 3711 4326 3741 4378
rect 3765 4326 3775 4378
rect 3775 4326 3821 4378
rect 3525 4324 3581 4326
rect 3605 4324 3661 4326
rect 3685 4324 3741 4326
rect 3765 4324 3821 4326
rect 3525 3290 3581 3292
rect 3605 3290 3661 3292
rect 3685 3290 3741 3292
rect 3765 3290 3821 3292
rect 3525 3238 3571 3290
rect 3571 3238 3581 3290
rect 3605 3238 3635 3290
rect 3635 3238 3647 3290
rect 3647 3238 3661 3290
rect 3685 3238 3699 3290
rect 3699 3238 3711 3290
rect 3711 3238 3741 3290
rect 3765 3238 3775 3290
rect 3775 3238 3821 3290
rect 3525 3236 3581 3238
rect 3605 3236 3661 3238
rect 3685 3236 3741 3238
rect 3765 3236 3821 3238
rect 7343 13082 7399 13084
rect 7423 13082 7479 13084
rect 7503 13082 7559 13084
rect 7583 13082 7639 13084
rect 7343 13030 7389 13082
rect 7389 13030 7399 13082
rect 7423 13030 7453 13082
rect 7453 13030 7465 13082
rect 7465 13030 7479 13082
rect 7503 13030 7517 13082
rect 7517 13030 7529 13082
rect 7529 13030 7559 13082
rect 7583 13030 7593 13082
rect 7593 13030 7639 13082
rect 7343 13028 7399 13030
rect 7423 13028 7479 13030
rect 7503 13028 7559 13030
rect 7583 13028 7639 13030
rect 10501 16890 10557 16892
rect 10581 16890 10637 16892
rect 10661 16890 10717 16892
rect 10741 16890 10797 16892
rect 10501 16838 10547 16890
rect 10547 16838 10557 16890
rect 10581 16838 10611 16890
rect 10611 16838 10623 16890
rect 10623 16838 10637 16890
rect 10661 16838 10675 16890
rect 10675 16838 10687 16890
rect 10687 16838 10717 16890
rect 10741 16838 10751 16890
rect 10751 16838 10797 16890
rect 10501 16836 10557 16838
rect 10581 16836 10637 16838
rect 10661 16836 10717 16838
rect 10741 16836 10797 16838
rect 11161 16346 11217 16348
rect 11241 16346 11297 16348
rect 11321 16346 11377 16348
rect 11401 16346 11457 16348
rect 11161 16294 11207 16346
rect 11207 16294 11217 16346
rect 11241 16294 11271 16346
rect 11271 16294 11283 16346
rect 11283 16294 11297 16346
rect 11321 16294 11335 16346
rect 11335 16294 11347 16346
rect 11347 16294 11377 16346
rect 11401 16294 11411 16346
rect 11411 16294 11457 16346
rect 11161 16292 11217 16294
rect 11241 16292 11297 16294
rect 11321 16292 11377 16294
rect 11401 16292 11457 16294
rect 14319 16890 14375 16892
rect 14399 16890 14455 16892
rect 14479 16890 14535 16892
rect 14559 16890 14615 16892
rect 14319 16838 14365 16890
rect 14365 16838 14375 16890
rect 14399 16838 14429 16890
rect 14429 16838 14441 16890
rect 14441 16838 14455 16890
rect 14479 16838 14493 16890
rect 14493 16838 14505 16890
rect 14505 16838 14535 16890
rect 14559 16838 14569 16890
rect 14569 16838 14615 16890
rect 14319 16836 14375 16838
rect 14399 16836 14455 16838
rect 14479 16836 14535 16838
rect 14559 16836 14615 16838
rect 10501 15802 10557 15804
rect 10581 15802 10637 15804
rect 10661 15802 10717 15804
rect 10741 15802 10797 15804
rect 10501 15750 10547 15802
rect 10547 15750 10557 15802
rect 10581 15750 10611 15802
rect 10611 15750 10623 15802
rect 10623 15750 10637 15802
rect 10661 15750 10675 15802
rect 10675 15750 10687 15802
rect 10687 15750 10717 15802
rect 10741 15750 10751 15802
rect 10751 15750 10797 15802
rect 10501 15748 10557 15750
rect 10581 15748 10637 15750
rect 10661 15748 10717 15750
rect 10741 15748 10797 15750
rect 11161 15258 11217 15260
rect 11241 15258 11297 15260
rect 11321 15258 11377 15260
rect 11401 15258 11457 15260
rect 11161 15206 11207 15258
rect 11207 15206 11217 15258
rect 11241 15206 11271 15258
rect 11271 15206 11283 15258
rect 11283 15206 11297 15258
rect 11321 15206 11335 15258
rect 11335 15206 11347 15258
rect 11347 15206 11377 15258
rect 11401 15206 11411 15258
rect 11411 15206 11457 15258
rect 11161 15204 11217 15206
rect 11241 15204 11297 15206
rect 11321 15204 11377 15206
rect 11401 15204 11457 15206
rect 14979 16346 15035 16348
rect 15059 16346 15115 16348
rect 15139 16346 15195 16348
rect 15219 16346 15275 16348
rect 14979 16294 15025 16346
rect 15025 16294 15035 16346
rect 15059 16294 15089 16346
rect 15089 16294 15101 16346
rect 15101 16294 15115 16346
rect 15139 16294 15153 16346
rect 15153 16294 15165 16346
rect 15165 16294 15195 16346
rect 15219 16294 15229 16346
rect 15229 16294 15275 16346
rect 14979 16292 15035 16294
rect 15059 16292 15115 16294
rect 15139 16292 15195 16294
rect 15219 16292 15275 16294
rect 10501 14714 10557 14716
rect 10581 14714 10637 14716
rect 10661 14714 10717 14716
rect 10741 14714 10797 14716
rect 10501 14662 10547 14714
rect 10547 14662 10557 14714
rect 10581 14662 10611 14714
rect 10611 14662 10623 14714
rect 10623 14662 10637 14714
rect 10661 14662 10675 14714
rect 10675 14662 10687 14714
rect 10687 14662 10717 14714
rect 10741 14662 10751 14714
rect 10751 14662 10797 14714
rect 10501 14660 10557 14662
rect 10581 14660 10637 14662
rect 10661 14660 10717 14662
rect 10741 14660 10797 14662
rect 6683 12538 6739 12540
rect 6763 12538 6819 12540
rect 6843 12538 6899 12540
rect 6923 12538 6979 12540
rect 6683 12486 6729 12538
rect 6729 12486 6739 12538
rect 6763 12486 6793 12538
rect 6793 12486 6805 12538
rect 6805 12486 6819 12538
rect 6843 12486 6857 12538
rect 6857 12486 6869 12538
rect 6869 12486 6899 12538
rect 6923 12486 6933 12538
rect 6933 12486 6979 12538
rect 6683 12484 6739 12486
rect 6763 12484 6819 12486
rect 6843 12484 6899 12486
rect 6923 12484 6979 12486
rect 6683 11450 6739 11452
rect 6763 11450 6819 11452
rect 6843 11450 6899 11452
rect 6923 11450 6979 11452
rect 6683 11398 6729 11450
rect 6729 11398 6739 11450
rect 6763 11398 6793 11450
rect 6793 11398 6805 11450
rect 6805 11398 6819 11450
rect 6843 11398 6857 11450
rect 6857 11398 6869 11450
rect 6869 11398 6899 11450
rect 6923 11398 6933 11450
rect 6933 11398 6979 11450
rect 6683 11396 6739 11398
rect 6763 11396 6819 11398
rect 6843 11396 6899 11398
rect 6923 11396 6979 11398
rect 7343 11994 7399 11996
rect 7423 11994 7479 11996
rect 7503 11994 7559 11996
rect 7583 11994 7639 11996
rect 7343 11942 7389 11994
rect 7389 11942 7399 11994
rect 7423 11942 7453 11994
rect 7453 11942 7465 11994
rect 7465 11942 7479 11994
rect 7503 11942 7517 11994
rect 7517 11942 7529 11994
rect 7529 11942 7559 11994
rect 7583 11942 7593 11994
rect 7593 11942 7639 11994
rect 7343 11940 7399 11942
rect 7423 11940 7479 11942
rect 7503 11940 7559 11942
rect 7583 11940 7639 11942
rect 7343 10906 7399 10908
rect 7423 10906 7479 10908
rect 7503 10906 7559 10908
rect 7583 10906 7639 10908
rect 7343 10854 7389 10906
rect 7389 10854 7399 10906
rect 7423 10854 7453 10906
rect 7453 10854 7465 10906
rect 7465 10854 7479 10906
rect 7503 10854 7517 10906
rect 7517 10854 7529 10906
rect 7529 10854 7559 10906
rect 7583 10854 7593 10906
rect 7593 10854 7639 10906
rect 7343 10852 7399 10854
rect 7423 10852 7479 10854
rect 7503 10852 7559 10854
rect 7583 10852 7639 10854
rect 6683 10362 6739 10364
rect 6763 10362 6819 10364
rect 6843 10362 6899 10364
rect 6923 10362 6979 10364
rect 6683 10310 6729 10362
rect 6729 10310 6739 10362
rect 6763 10310 6793 10362
rect 6793 10310 6805 10362
rect 6805 10310 6819 10362
rect 6843 10310 6857 10362
rect 6857 10310 6869 10362
rect 6869 10310 6899 10362
rect 6923 10310 6933 10362
rect 6933 10310 6979 10362
rect 6683 10308 6739 10310
rect 6763 10308 6819 10310
rect 6843 10308 6899 10310
rect 6923 10308 6979 10310
rect 5446 7248 5502 7304
rect 6683 9274 6739 9276
rect 6763 9274 6819 9276
rect 6843 9274 6899 9276
rect 6923 9274 6979 9276
rect 6683 9222 6729 9274
rect 6729 9222 6739 9274
rect 6763 9222 6793 9274
rect 6793 9222 6805 9274
rect 6805 9222 6819 9274
rect 6843 9222 6857 9274
rect 6857 9222 6869 9274
rect 6869 9222 6899 9274
rect 6923 9222 6933 9274
rect 6933 9222 6979 9274
rect 6683 9220 6739 9222
rect 6763 9220 6819 9222
rect 6843 9220 6899 9222
rect 6923 9220 6979 9222
rect 6683 8186 6739 8188
rect 6763 8186 6819 8188
rect 6843 8186 6899 8188
rect 6923 8186 6979 8188
rect 6683 8134 6729 8186
rect 6729 8134 6739 8186
rect 6763 8134 6793 8186
rect 6793 8134 6805 8186
rect 6805 8134 6819 8186
rect 6843 8134 6857 8186
rect 6857 8134 6869 8186
rect 6869 8134 6899 8186
rect 6923 8134 6933 8186
rect 6933 8134 6979 8186
rect 6683 8132 6739 8134
rect 6763 8132 6819 8134
rect 6843 8132 6899 8134
rect 6923 8132 6979 8134
rect 6683 7098 6739 7100
rect 6763 7098 6819 7100
rect 6843 7098 6899 7100
rect 6923 7098 6979 7100
rect 6683 7046 6729 7098
rect 6729 7046 6739 7098
rect 6763 7046 6793 7098
rect 6793 7046 6805 7098
rect 6805 7046 6819 7098
rect 6843 7046 6857 7098
rect 6857 7046 6869 7098
rect 6869 7046 6899 7098
rect 6923 7046 6933 7098
rect 6933 7046 6979 7098
rect 6683 7044 6739 7046
rect 6763 7044 6819 7046
rect 6843 7044 6899 7046
rect 6923 7044 6979 7046
rect 7343 9818 7399 9820
rect 7423 9818 7479 9820
rect 7503 9818 7559 9820
rect 7583 9818 7639 9820
rect 7343 9766 7389 9818
rect 7389 9766 7399 9818
rect 7423 9766 7453 9818
rect 7453 9766 7465 9818
rect 7465 9766 7479 9818
rect 7503 9766 7517 9818
rect 7517 9766 7529 9818
rect 7529 9766 7559 9818
rect 7583 9766 7593 9818
rect 7593 9766 7639 9818
rect 7343 9764 7399 9766
rect 7423 9764 7479 9766
rect 7503 9764 7559 9766
rect 7583 9764 7639 9766
rect 7470 9560 7526 9616
rect 7470 9052 7472 9072
rect 7472 9052 7524 9072
rect 7524 9052 7526 9072
rect 7470 9016 7526 9052
rect 7343 8730 7399 8732
rect 7423 8730 7479 8732
rect 7503 8730 7559 8732
rect 7583 8730 7639 8732
rect 7343 8678 7389 8730
rect 7389 8678 7399 8730
rect 7423 8678 7453 8730
rect 7453 8678 7465 8730
rect 7465 8678 7479 8730
rect 7503 8678 7517 8730
rect 7517 8678 7529 8730
rect 7529 8678 7559 8730
rect 7583 8678 7593 8730
rect 7593 8678 7639 8730
rect 7343 8676 7399 8678
rect 7423 8676 7479 8678
rect 7503 8676 7559 8678
rect 7583 8676 7639 8678
rect 6683 6010 6739 6012
rect 6763 6010 6819 6012
rect 6843 6010 6899 6012
rect 6923 6010 6979 6012
rect 6683 5958 6729 6010
rect 6729 5958 6739 6010
rect 6763 5958 6793 6010
rect 6793 5958 6805 6010
rect 6805 5958 6819 6010
rect 6843 5958 6857 6010
rect 6857 5958 6869 6010
rect 6869 5958 6899 6010
rect 6923 5958 6933 6010
rect 6933 5958 6979 6010
rect 6683 5956 6739 5958
rect 6763 5956 6819 5958
rect 6843 5956 6899 5958
rect 6923 5956 6979 5958
rect 6683 4922 6739 4924
rect 6763 4922 6819 4924
rect 6843 4922 6899 4924
rect 6923 4922 6979 4924
rect 6683 4870 6729 4922
rect 6729 4870 6739 4922
rect 6763 4870 6793 4922
rect 6793 4870 6805 4922
rect 6805 4870 6819 4922
rect 6843 4870 6857 4922
rect 6857 4870 6869 4922
rect 6869 4870 6899 4922
rect 6923 4870 6933 4922
rect 6933 4870 6979 4922
rect 6683 4868 6739 4870
rect 6763 4868 6819 4870
rect 6843 4868 6899 4870
rect 6923 4868 6979 4870
rect 7343 7642 7399 7644
rect 7423 7642 7479 7644
rect 7503 7642 7559 7644
rect 7583 7642 7639 7644
rect 7343 7590 7389 7642
rect 7389 7590 7399 7642
rect 7423 7590 7453 7642
rect 7453 7590 7465 7642
rect 7465 7590 7479 7642
rect 7503 7590 7517 7642
rect 7517 7590 7529 7642
rect 7529 7590 7559 7642
rect 7583 7590 7593 7642
rect 7593 7590 7639 7642
rect 7343 7588 7399 7590
rect 7423 7588 7479 7590
rect 7503 7588 7559 7590
rect 7583 7588 7639 7590
rect 10501 13626 10557 13628
rect 10581 13626 10637 13628
rect 10661 13626 10717 13628
rect 10741 13626 10797 13628
rect 10501 13574 10547 13626
rect 10547 13574 10557 13626
rect 10581 13574 10611 13626
rect 10611 13574 10623 13626
rect 10623 13574 10637 13626
rect 10661 13574 10675 13626
rect 10675 13574 10687 13626
rect 10687 13574 10717 13626
rect 10741 13574 10751 13626
rect 10751 13574 10797 13626
rect 10501 13572 10557 13574
rect 10581 13572 10637 13574
rect 10661 13572 10717 13574
rect 10741 13572 10797 13574
rect 11161 14170 11217 14172
rect 11241 14170 11297 14172
rect 11321 14170 11377 14172
rect 11401 14170 11457 14172
rect 11161 14118 11207 14170
rect 11207 14118 11217 14170
rect 11241 14118 11271 14170
rect 11271 14118 11283 14170
rect 11283 14118 11297 14170
rect 11321 14118 11335 14170
rect 11335 14118 11347 14170
rect 11347 14118 11377 14170
rect 11401 14118 11411 14170
rect 11411 14118 11457 14170
rect 11161 14116 11217 14118
rect 11241 14116 11297 14118
rect 11321 14116 11377 14118
rect 11401 14116 11457 14118
rect 11161 13082 11217 13084
rect 11241 13082 11297 13084
rect 11321 13082 11377 13084
rect 11401 13082 11457 13084
rect 11161 13030 11207 13082
rect 11207 13030 11217 13082
rect 11241 13030 11271 13082
rect 11271 13030 11283 13082
rect 11283 13030 11297 13082
rect 11321 13030 11335 13082
rect 11335 13030 11347 13082
rect 11347 13030 11377 13082
rect 11401 13030 11411 13082
rect 11411 13030 11457 13082
rect 11161 13028 11217 13030
rect 11241 13028 11297 13030
rect 11321 13028 11377 13030
rect 11401 13028 11457 13030
rect 10501 12538 10557 12540
rect 10581 12538 10637 12540
rect 10661 12538 10717 12540
rect 10741 12538 10797 12540
rect 10501 12486 10547 12538
rect 10547 12486 10557 12538
rect 10581 12486 10611 12538
rect 10611 12486 10623 12538
rect 10623 12486 10637 12538
rect 10661 12486 10675 12538
rect 10675 12486 10687 12538
rect 10687 12486 10717 12538
rect 10741 12486 10751 12538
rect 10751 12486 10797 12538
rect 10501 12484 10557 12486
rect 10581 12484 10637 12486
rect 10661 12484 10717 12486
rect 10741 12484 10797 12486
rect 11161 11994 11217 11996
rect 11241 11994 11297 11996
rect 11321 11994 11377 11996
rect 11401 11994 11457 11996
rect 11161 11942 11207 11994
rect 11207 11942 11217 11994
rect 11241 11942 11271 11994
rect 11271 11942 11283 11994
rect 11283 11942 11297 11994
rect 11321 11942 11335 11994
rect 11335 11942 11347 11994
rect 11347 11942 11377 11994
rect 11401 11942 11411 11994
rect 11411 11942 11457 11994
rect 11161 11940 11217 11942
rect 11241 11940 11297 11942
rect 11321 11940 11377 11942
rect 11401 11940 11457 11942
rect 14319 15802 14375 15804
rect 14399 15802 14455 15804
rect 14479 15802 14535 15804
rect 14559 15802 14615 15804
rect 14319 15750 14365 15802
rect 14365 15750 14375 15802
rect 14399 15750 14429 15802
rect 14429 15750 14441 15802
rect 14441 15750 14455 15802
rect 14479 15750 14493 15802
rect 14493 15750 14505 15802
rect 14505 15750 14535 15802
rect 14559 15750 14569 15802
rect 14569 15750 14615 15802
rect 14319 15748 14375 15750
rect 14399 15748 14455 15750
rect 14479 15748 14535 15750
rect 14559 15748 14615 15750
rect 14979 15258 15035 15260
rect 15059 15258 15115 15260
rect 15139 15258 15195 15260
rect 15219 15258 15275 15260
rect 14979 15206 15025 15258
rect 15025 15206 15035 15258
rect 15059 15206 15089 15258
rect 15089 15206 15101 15258
rect 15101 15206 15115 15258
rect 15139 15206 15153 15258
rect 15153 15206 15165 15258
rect 15165 15206 15195 15258
rect 15219 15206 15229 15258
rect 15229 15206 15275 15258
rect 14979 15204 15035 15206
rect 15059 15204 15115 15206
rect 15139 15204 15195 15206
rect 15219 15204 15275 15206
rect 16026 15000 16082 15056
rect 14319 14714 14375 14716
rect 14399 14714 14455 14716
rect 14479 14714 14535 14716
rect 14559 14714 14615 14716
rect 14319 14662 14365 14714
rect 14365 14662 14375 14714
rect 14399 14662 14429 14714
rect 14429 14662 14441 14714
rect 14441 14662 14455 14714
rect 14479 14662 14493 14714
rect 14493 14662 14505 14714
rect 14505 14662 14535 14714
rect 14559 14662 14569 14714
rect 14569 14662 14615 14714
rect 14319 14660 14375 14662
rect 14399 14660 14455 14662
rect 14479 14660 14535 14662
rect 14559 14660 14615 14662
rect 14979 14170 15035 14172
rect 15059 14170 15115 14172
rect 15139 14170 15195 14172
rect 15219 14170 15275 14172
rect 14979 14118 15025 14170
rect 15025 14118 15035 14170
rect 15059 14118 15089 14170
rect 15089 14118 15101 14170
rect 15101 14118 15115 14170
rect 15139 14118 15153 14170
rect 15153 14118 15165 14170
rect 15165 14118 15195 14170
rect 15219 14118 15229 14170
rect 15229 14118 15275 14170
rect 14979 14116 15035 14118
rect 15059 14116 15115 14118
rect 15139 14116 15195 14118
rect 15219 14116 15275 14118
rect 14319 13626 14375 13628
rect 14399 13626 14455 13628
rect 14479 13626 14535 13628
rect 14559 13626 14615 13628
rect 14319 13574 14365 13626
rect 14365 13574 14375 13626
rect 14399 13574 14429 13626
rect 14429 13574 14441 13626
rect 14441 13574 14455 13626
rect 14479 13574 14493 13626
rect 14493 13574 14505 13626
rect 14505 13574 14535 13626
rect 14559 13574 14569 13626
rect 14569 13574 14615 13626
rect 14319 13572 14375 13574
rect 14399 13572 14455 13574
rect 14479 13572 14535 13574
rect 14559 13572 14615 13574
rect 14979 13082 15035 13084
rect 15059 13082 15115 13084
rect 15139 13082 15195 13084
rect 15219 13082 15275 13084
rect 14979 13030 15025 13082
rect 15025 13030 15035 13082
rect 15059 13030 15089 13082
rect 15089 13030 15101 13082
rect 15101 13030 15115 13082
rect 15139 13030 15153 13082
rect 15153 13030 15165 13082
rect 15165 13030 15195 13082
rect 15219 13030 15229 13082
rect 15229 13030 15275 13082
rect 14979 13028 15035 13030
rect 15059 13028 15115 13030
rect 15139 13028 15195 13030
rect 15219 13028 15275 13030
rect 15934 12960 15990 13016
rect 14319 12538 14375 12540
rect 14399 12538 14455 12540
rect 14479 12538 14535 12540
rect 14559 12538 14615 12540
rect 14319 12486 14365 12538
rect 14365 12486 14375 12538
rect 14399 12486 14429 12538
rect 14429 12486 14441 12538
rect 14441 12486 14455 12538
rect 14479 12486 14493 12538
rect 14493 12486 14505 12538
rect 14505 12486 14535 12538
rect 14559 12486 14569 12538
rect 14569 12486 14615 12538
rect 14319 12484 14375 12486
rect 14399 12484 14455 12486
rect 14479 12484 14535 12486
rect 14559 12484 14615 12486
rect 10501 11450 10557 11452
rect 10581 11450 10637 11452
rect 10661 11450 10717 11452
rect 10741 11450 10797 11452
rect 10501 11398 10547 11450
rect 10547 11398 10557 11450
rect 10581 11398 10611 11450
rect 10611 11398 10623 11450
rect 10623 11398 10637 11450
rect 10661 11398 10675 11450
rect 10675 11398 10687 11450
rect 10687 11398 10717 11450
rect 10741 11398 10751 11450
rect 10751 11398 10797 11450
rect 10501 11396 10557 11398
rect 10581 11396 10637 11398
rect 10661 11396 10717 11398
rect 10741 11396 10797 11398
rect 8390 9052 8392 9072
rect 8392 9052 8444 9072
rect 8444 9052 8446 9072
rect 8390 9016 8446 9052
rect 11161 10906 11217 10908
rect 11241 10906 11297 10908
rect 11321 10906 11377 10908
rect 11401 10906 11457 10908
rect 11161 10854 11207 10906
rect 11207 10854 11217 10906
rect 11241 10854 11271 10906
rect 11271 10854 11283 10906
rect 11283 10854 11297 10906
rect 11321 10854 11335 10906
rect 11335 10854 11347 10906
rect 11347 10854 11377 10906
rect 11401 10854 11411 10906
rect 11411 10854 11457 10906
rect 11161 10852 11217 10854
rect 11241 10852 11297 10854
rect 11321 10852 11377 10854
rect 11401 10852 11457 10854
rect 10501 10362 10557 10364
rect 10581 10362 10637 10364
rect 10661 10362 10717 10364
rect 10741 10362 10797 10364
rect 10501 10310 10547 10362
rect 10547 10310 10557 10362
rect 10581 10310 10611 10362
rect 10611 10310 10623 10362
rect 10623 10310 10637 10362
rect 10661 10310 10675 10362
rect 10675 10310 10687 10362
rect 10687 10310 10717 10362
rect 10741 10310 10751 10362
rect 10751 10310 10797 10362
rect 10501 10308 10557 10310
rect 10581 10308 10637 10310
rect 10661 10308 10717 10310
rect 10741 10308 10797 10310
rect 14979 11994 15035 11996
rect 15059 11994 15115 11996
rect 15139 11994 15195 11996
rect 15219 11994 15275 11996
rect 14979 11942 15025 11994
rect 15025 11942 15035 11994
rect 15059 11942 15089 11994
rect 15089 11942 15101 11994
rect 15101 11942 15115 11994
rect 15139 11942 15153 11994
rect 15153 11942 15165 11994
rect 15165 11942 15195 11994
rect 15219 11942 15229 11994
rect 15229 11942 15275 11994
rect 14979 11940 15035 11942
rect 15059 11940 15115 11942
rect 15139 11940 15195 11942
rect 15219 11940 15275 11942
rect 9034 9596 9036 9616
rect 9036 9596 9088 9616
rect 9088 9596 9090 9616
rect 9034 9560 9090 9596
rect 7343 6554 7399 6556
rect 7423 6554 7479 6556
rect 7503 6554 7559 6556
rect 7583 6554 7639 6556
rect 7343 6502 7389 6554
rect 7389 6502 7399 6554
rect 7423 6502 7453 6554
rect 7453 6502 7465 6554
rect 7465 6502 7479 6554
rect 7503 6502 7517 6554
rect 7517 6502 7529 6554
rect 7529 6502 7559 6554
rect 7583 6502 7593 6554
rect 7593 6502 7639 6554
rect 7343 6500 7399 6502
rect 7423 6500 7479 6502
rect 7503 6500 7559 6502
rect 7583 6500 7639 6502
rect 7343 5466 7399 5468
rect 7423 5466 7479 5468
rect 7503 5466 7559 5468
rect 7583 5466 7639 5468
rect 7343 5414 7389 5466
rect 7389 5414 7399 5466
rect 7423 5414 7453 5466
rect 7453 5414 7465 5466
rect 7465 5414 7479 5466
rect 7503 5414 7517 5466
rect 7517 5414 7529 5466
rect 7529 5414 7559 5466
rect 7583 5414 7593 5466
rect 7593 5414 7639 5466
rect 7343 5412 7399 5414
rect 7423 5412 7479 5414
rect 7503 5412 7559 5414
rect 7583 5412 7639 5414
rect 6683 3834 6739 3836
rect 6763 3834 6819 3836
rect 6843 3834 6899 3836
rect 6923 3834 6979 3836
rect 6683 3782 6729 3834
rect 6729 3782 6739 3834
rect 6763 3782 6793 3834
rect 6793 3782 6805 3834
rect 6805 3782 6819 3834
rect 6843 3782 6857 3834
rect 6857 3782 6869 3834
rect 6869 3782 6899 3834
rect 6923 3782 6933 3834
rect 6933 3782 6979 3834
rect 6683 3780 6739 3782
rect 6763 3780 6819 3782
rect 6843 3780 6899 3782
rect 6923 3780 6979 3782
rect 6090 3596 6146 3632
rect 6090 3576 6092 3596
rect 6092 3576 6144 3596
rect 6144 3576 6146 3596
rect 6734 3612 6736 3632
rect 6736 3612 6788 3632
rect 6788 3612 6790 3632
rect 6734 3576 6790 3612
rect 938 2760 994 2816
rect 2865 2746 2921 2748
rect 2945 2746 3001 2748
rect 3025 2746 3081 2748
rect 3105 2746 3161 2748
rect 2865 2694 2911 2746
rect 2911 2694 2921 2746
rect 2945 2694 2975 2746
rect 2975 2694 2987 2746
rect 2987 2694 3001 2746
rect 3025 2694 3039 2746
rect 3039 2694 3051 2746
rect 3051 2694 3081 2746
rect 3105 2694 3115 2746
rect 3115 2694 3161 2746
rect 2865 2692 2921 2694
rect 2945 2692 3001 2694
rect 3025 2692 3081 2694
rect 3105 2692 3161 2694
rect 6683 2746 6739 2748
rect 6763 2746 6819 2748
rect 6843 2746 6899 2748
rect 6923 2746 6979 2748
rect 6683 2694 6729 2746
rect 6729 2694 6739 2746
rect 6763 2694 6793 2746
rect 6793 2694 6805 2746
rect 6805 2694 6819 2746
rect 6843 2694 6857 2746
rect 6857 2694 6869 2746
rect 6869 2694 6899 2746
rect 6923 2694 6933 2746
rect 6933 2694 6979 2746
rect 6683 2692 6739 2694
rect 6763 2692 6819 2694
rect 6843 2692 6899 2694
rect 6923 2692 6979 2694
rect 7343 4378 7399 4380
rect 7423 4378 7479 4380
rect 7503 4378 7559 4380
rect 7583 4378 7639 4380
rect 7343 4326 7389 4378
rect 7389 4326 7399 4378
rect 7423 4326 7453 4378
rect 7453 4326 7465 4378
rect 7465 4326 7479 4378
rect 7503 4326 7517 4378
rect 7517 4326 7529 4378
rect 7529 4326 7559 4378
rect 7583 4326 7593 4378
rect 7593 4326 7639 4378
rect 7343 4324 7399 4326
rect 7423 4324 7479 4326
rect 7503 4324 7559 4326
rect 7583 4324 7639 4326
rect 7343 3290 7399 3292
rect 7423 3290 7479 3292
rect 7503 3290 7559 3292
rect 7583 3290 7639 3292
rect 7343 3238 7389 3290
rect 7389 3238 7399 3290
rect 7423 3238 7453 3290
rect 7453 3238 7465 3290
rect 7465 3238 7479 3290
rect 7503 3238 7517 3290
rect 7517 3238 7529 3290
rect 7529 3238 7559 3290
rect 7583 3238 7593 3290
rect 7593 3238 7639 3290
rect 7343 3236 7399 3238
rect 7423 3236 7479 3238
rect 7503 3236 7559 3238
rect 7583 3236 7639 3238
rect 11161 9818 11217 9820
rect 11241 9818 11297 9820
rect 11321 9818 11377 9820
rect 11401 9818 11457 9820
rect 11161 9766 11207 9818
rect 11207 9766 11217 9818
rect 11241 9766 11271 9818
rect 11271 9766 11283 9818
rect 11283 9766 11297 9818
rect 11321 9766 11335 9818
rect 11335 9766 11347 9818
rect 11347 9766 11377 9818
rect 11401 9766 11411 9818
rect 11411 9766 11457 9818
rect 11161 9764 11217 9766
rect 11241 9764 11297 9766
rect 11321 9764 11377 9766
rect 11401 9764 11457 9766
rect 10501 9274 10557 9276
rect 10581 9274 10637 9276
rect 10661 9274 10717 9276
rect 10741 9274 10797 9276
rect 10501 9222 10547 9274
rect 10547 9222 10557 9274
rect 10581 9222 10611 9274
rect 10611 9222 10623 9274
rect 10623 9222 10637 9274
rect 10661 9222 10675 9274
rect 10675 9222 10687 9274
rect 10687 9222 10717 9274
rect 10741 9222 10751 9274
rect 10751 9222 10797 9274
rect 10501 9220 10557 9222
rect 10581 9220 10637 9222
rect 10661 9220 10717 9222
rect 10741 9220 10797 9222
rect 11161 8730 11217 8732
rect 11241 8730 11297 8732
rect 11321 8730 11377 8732
rect 11401 8730 11457 8732
rect 11161 8678 11207 8730
rect 11207 8678 11217 8730
rect 11241 8678 11271 8730
rect 11271 8678 11283 8730
rect 11283 8678 11297 8730
rect 11321 8678 11335 8730
rect 11335 8678 11347 8730
rect 11347 8678 11377 8730
rect 11401 8678 11411 8730
rect 11411 8678 11457 8730
rect 11161 8676 11217 8678
rect 11241 8676 11297 8678
rect 11321 8676 11377 8678
rect 11401 8676 11457 8678
rect 10501 8186 10557 8188
rect 10581 8186 10637 8188
rect 10661 8186 10717 8188
rect 10741 8186 10797 8188
rect 10501 8134 10547 8186
rect 10547 8134 10557 8186
rect 10581 8134 10611 8186
rect 10611 8134 10623 8186
rect 10623 8134 10637 8186
rect 10661 8134 10675 8186
rect 10675 8134 10687 8186
rect 10687 8134 10717 8186
rect 10741 8134 10751 8186
rect 10751 8134 10797 8186
rect 10501 8132 10557 8134
rect 10581 8132 10637 8134
rect 10661 8132 10717 8134
rect 10741 8132 10797 8134
rect 11161 7642 11217 7644
rect 11241 7642 11297 7644
rect 11321 7642 11377 7644
rect 11401 7642 11457 7644
rect 11161 7590 11207 7642
rect 11207 7590 11217 7642
rect 11241 7590 11271 7642
rect 11271 7590 11283 7642
rect 11283 7590 11297 7642
rect 11321 7590 11335 7642
rect 11335 7590 11347 7642
rect 11347 7590 11377 7642
rect 11401 7590 11411 7642
rect 11411 7590 11457 7642
rect 11161 7588 11217 7590
rect 11241 7588 11297 7590
rect 11321 7588 11377 7590
rect 11401 7588 11457 7590
rect 10501 7098 10557 7100
rect 10581 7098 10637 7100
rect 10661 7098 10717 7100
rect 10741 7098 10797 7100
rect 10501 7046 10547 7098
rect 10547 7046 10557 7098
rect 10581 7046 10611 7098
rect 10611 7046 10623 7098
rect 10623 7046 10637 7098
rect 10661 7046 10675 7098
rect 10675 7046 10687 7098
rect 10687 7046 10717 7098
rect 10741 7046 10751 7098
rect 10751 7046 10797 7098
rect 10501 7044 10557 7046
rect 10581 7044 10637 7046
rect 10661 7044 10717 7046
rect 10741 7044 10797 7046
rect 14319 11450 14375 11452
rect 14399 11450 14455 11452
rect 14479 11450 14535 11452
rect 14559 11450 14615 11452
rect 14319 11398 14365 11450
rect 14365 11398 14375 11450
rect 14399 11398 14429 11450
rect 14429 11398 14441 11450
rect 14441 11398 14455 11450
rect 14479 11398 14493 11450
rect 14493 11398 14505 11450
rect 14505 11398 14535 11450
rect 14559 11398 14569 11450
rect 14569 11398 14615 11450
rect 14319 11396 14375 11398
rect 14399 11396 14455 11398
rect 14479 11396 14535 11398
rect 14559 11396 14615 11398
rect 11161 6554 11217 6556
rect 11241 6554 11297 6556
rect 11321 6554 11377 6556
rect 11401 6554 11457 6556
rect 11161 6502 11207 6554
rect 11207 6502 11217 6554
rect 11241 6502 11271 6554
rect 11271 6502 11283 6554
rect 11283 6502 11297 6554
rect 11321 6502 11335 6554
rect 11335 6502 11347 6554
rect 11347 6502 11377 6554
rect 11401 6502 11411 6554
rect 11411 6502 11457 6554
rect 11161 6500 11217 6502
rect 11241 6500 11297 6502
rect 11321 6500 11377 6502
rect 11401 6500 11457 6502
rect 14319 10362 14375 10364
rect 14399 10362 14455 10364
rect 14479 10362 14535 10364
rect 14559 10362 14615 10364
rect 14319 10310 14365 10362
rect 14365 10310 14375 10362
rect 14399 10310 14429 10362
rect 14429 10310 14441 10362
rect 14441 10310 14455 10362
rect 14479 10310 14493 10362
rect 14493 10310 14505 10362
rect 14505 10310 14535 10362
rect 14559 10310 14569 10362
rect 14569 10310 14615 10362
rect 14319 10308 14375 10310
rect 14399 10308 14455 10310
rect 14479 10308 14535 10310
rect 14559 10308 14615 10310
rect 14979 10906 15035 10908
rect 15059 10906 15115 10908
rect 15139 10906 15195 10908
rect 15219 10906 15275 10908
rect 14979 10854 15025 10906
rect 15025 10854 15035 10906
rect 15059 10854 15089 10906
rect 15089 10854 15101 10906
rect 15101 10854 15115 10906
rect 15139 10854 15153 10906
rect 15153 10854 15165 10906
rect 15165 10854 15195 10906
rect 15219 10854 15229 10906
rect 15229 10854 15275 10906
rect 14979 10852 15035 10854
rect 15059 10852 15115 10854
rect 15139 10852 15195 10854
rect 15219 10852 15275 10854
rect 16026 10920 16082 10976
rect 14319 9274 14375 9276
rect 14399 9274 14455 9276
rect 14479 9274 14535 9276
rect 14559 9274 14615 9276
rect 14319 9222 14365 9274
rect 14365 9222 14375 9274
rect 14399 9222 14429 9274
rect 14429 9222 14441 9274
rect 14441 9222 14455 9274
rect 14479 9222 14493 9274
rect 14493 9222 14505 9274
rect 14505 9222 14535 9274
rect 14559 9222 14569 9274
rect 14569 9222 14615 9274
rect 14319 9220 14375 9222
rect 14399 9220 14455 9222
rect 14479 9220 14535 9222
rect 14559 9220 14615 9222
rect 14979 9818 15035 9820
rect 15059 9818 15115 9820
rect 15139 9818 15195 9820
rect 15219 9818 15275 9820
rect 14979 9766 15025 9818
rect 15025 9766 15035 9818
rect 15059 9766 15089 9818
rect 15089 9766 15101 9818
rect 15101 9766 15115 9818
rect 15139 9766 15153 9818
rect 15153 9766 15165 9818
rect 15165 9766 15195 9818
rect 15219 9766 15229 9818
rect 15229 9766 15275 9818
rect 14979 9764 15035 9766
rect 15059 9764 15115 9766
rect 15139 9764 15195 9766
rect 15219 9764 15275 9766
rect 14979 8730 15035 8732
rect 15059 8730 15115 8732
rect 15139 8730 15195 8732
rect 15219 8730 15275 8732
rect 14979 8678 15025 8730
rect 15025 8678 15035 8730
rect 15059 8678 15089 8730
rect 15089 8678 15101 8730
rect 15101 8678 15115 8730
rect 15139 8678 15153 8730
rect 15153 8678 15165 8730
rect 15165 8678 15195 8730
rect 15219 8678 15229 8730
rect 15229 8678 15275 8730
rect 14979 8676 15035 8678
rect 15059 8676 15115 8678
rect 15139 8676 15195 8678
rect 15219 8676 15275 8678
rect 16026 9560 16082 9616
rect 14319 8186 14375 8188
rect 14399 8186 14455 8188
rect 14479 8186 14535 8188
rect 14559 8186 14615 8188
rect 14319 8134 14365 8186
rect 14365 8134 14375 8186
rect 14399 8134 14429 8186
rect 14429 8134 14441 8186
rect 14441 8134 14455 8186
rect 14479 8134 14493 8186
rect 14493 8134 14505 8186
rect 14505 8134 14535 8186
rect 14559 8134 14569 8186
rect 14569 8134 14615 8186
rect 14319 8132 14375 8134
rect 14399 8132 14455 8134
rect 14479 8132 14535 8134
rect 14559 8132 14615 8134
rect 14319 7098 14375 7100
rect 14399 7098 14455 7100
rect 14479 7098 14535 7100
rect 14559 7098 14615 7100
rect 14319 7046 14365 7098
rect 14365 7046 14375 7098
rect 14399 7046 14429 7098
rect 14429 7046 14441 7098
rect 14441 7046 14455 7098
rect 14479 7046 14493 7098
rect 14493 7046 14505 7098
rect 14505 7046 14535 7098
rect 14559 7046 14569 7098
rect 14569 7046 14615 7098
rect 14319 7044 14375 7046
rect 14399 7044 14455 7046
rect 14479 7044 14535 7046
rect 14559 7044 14615 7046
rect 14979 7642 15035 7644
rect 15059 7642 15115 7644
rect 15139 7642 15195 7644
rect 15219 7642 15275 7644
rect 14979 7590 15025 7642
rect 15025 7590 15035 7642
rect 15059 7590 15089 7642
rect 15089 7590 15101 7642
rect 15101 7590 15115 7642
rect 15139 7590 15153 7642
rect 15153 7590 15165 7642
rect 15165 7590 15195 7642
rect 15219 7590 15229 7642
rect 15229 7590 15275 7642
rect 14979 7588 15035 7590
rect 15059 7588 15115 7590
rect 15139 7588 15195 7590
rect 15219 7588 15275 7590
rect 15934 7520 15990 7576
rect 14979 6554 15035 6556
rect 15059 6554 15115 6556
rect 15139 6554 15195 6556
rect 15219 6554 15275 6556
rect 14979 6502 15025 6554
rect 15025 6502 15035 6554
rect 15059 6502 15089 6554
rect 15089 6502 15101 6554
rect 15101 6502 15115 6554
rect 15139 6502 15153 6554
rect 15153 6502 15165 6554
rect 15165 6502 15195 6554
rect 15219 6502 15229 6554
rect 15229 6502 15275 6554
rect 14979 6500 15035 6502
rect 15059 6500 15115 6502
rect 15139 6500 15195 6502
rect 15219 6500 15275 6502
rect 10501 6010 10557 6012
rect 10581 6010 10637 6012
rect 10661 6010 10717 6012
rect 10741 6010 10797 6012
rect 10501 5958 10547 6010
rect 10547 5958 10557 6010
rect 10581 5958 10611 6010
rect 10611 5958 10623 6010
rect 10623 5958 10637 6010
rect 10661 5958 10675 6010
rect 10675 5958 10687 6010
rect 10687 5958 10717 6010
rect 10741 5958 10751 6010
rect 10751 5958 10797 6010
rect 10501 5956 10557 5958
rect 10581 5956 10637 5958
rect 10661 5956 10717 5958
rect 10741 5956 10797 5958
rect 11161 5466 11217 5468
rect 11241 5466 11297 5468
rect 11321 5466 11377 5468
rect 11401 5466 11457 5468
rect 11161 5414 11207 5466
rect 11207 5414 11217 5466
rect 11241 5414 11271 5466
rect 11271 5414 11283 5466
rect 11283 5414 11297 5466
rect 11321 5414 11335 5466
rect 11335 5414 11347 5466
rect 11347 5414 11377 5466
rect 11401 5414 11411 5466
rect 11411 5414 11457 5466
rect 11161 5412 11217 5414
rect 11241 5412 11297 5414
rect 11321 5412 11377 5414
rect 11401 5412 11457 5414
rect 10501 4922 10557 4924
rect 10581 4922 10637 4924
rect 10661 4922 10717 4924
rect 10741 4922 10797 4924
rect 10501 4870 10547 4922
rect 10547 4870 10557 4922
rect 10581 4870 10611 4922
rect 10611 4870 10623 4922
rect 10623 4870 10637 4922
rect 10661 4870 10675 4922
rect 10675 4870 10687 4922
rect 10687 4870 10717 4922
rect 10741 4870 10751 4922
rect 10751 4870 10797 4922
rect 10501 4868 10557 4870
rect 10581 4868 10637 4870
rect 10661 4868 10717 4870
rect 10741 4868 10797 4870
rect 11161 4378 11217 4380
rect 11241 4378 11297 4380
rect 11321 4378 11377 4380
rect 11401 4378 11457 4380
rect 11161 4326 11207 4378
rect 11207 4326 11217 4378
rect 11241 4326 11271 4378
rect 11271 4326 11283 4378
rect 11283 4326 11297 4378
rect 11321 4326 11335 4378
rect 11335 4326 11347 4378
rect 11347 4326 11377 4378
rect 11401 4326 11411 4378
rect 11411 4326 11457 4378
rect 11161 4324 11217 4326
rect 11241 4324 11297 4326
rect 11321 4324 11377 4326
rect 11401 4324 11457 4326
rect 14319 6010 14375 6012
rect 14399 6010 14455 6012
rect 14479 6010 14535 6012
rect 14559 6010 14615 6012
rect 14319 5958 14365 6010
rect 14365 5958 14375 6010
rect 14399 5958 14429 6010
rect 14429 5958 14441 6010
rect 14441 5958 14455 6010
rect 14479 5958 14493 6010
rect 14493 5958 14505 6010
rect 14505 5958 14535 6010
rect 14559 5958 14569 6010
rect 14569 5958 14615 6010
rect 14319 5956 14375 5958
rect 14399 5956 14455 5958
rect 14479 5956 14535 5958
rect 14559 5956 14615 5958
rect 14319 4922 14375 4924
rect 14399 4922 14455 4924
rect 14479 4922 14535 4924
rect 14559 4922 14615 4924
rect 14319 4870 14365 4922
rect 14365 4870 14375 4922
rect 14399 4870 14429 4922
rect 14429 4870 14441 4922
rect 14441 4870 14455 4922
rect 14479 4870 14493 4922
rect 14493 4870 14505 4922
rect 14505 4870 14535 4922
rect 14559 4870 14569 4922
rect 14569 4870 14615 4922
rect 14319 4868 14375 4870
rect 14399 4868 14455 4870
rect 14479 4868 14535 4870
rect 14559 4868 14615 4870
rect 16026 5516 16028 5536
rect 16028 5516 16080 5536
rect 16080 5516 16082 5536
rect 16026 5480 16082 5516
rect 14979 5466 15035 5468
rect 15059 5466 15115 5468
rect 15139 5466 15195 5468
rect 15219 5466 15275 5468
rect 14979 5414 15025 5466
rect 15025 5414 15035 5466
rect 15059 5414 15089 5466
rect 15089 5414 15101 5466
rect 15101 5414 15115 5466
rect 15139 5414 15153 5466
rect 15153 5414 15165 5466
rect 15165 5414 15195 5466
rect 15219 5414 15229 5466
rect 15229 5414 15275 5466
rect 14979 5412 15035 5414
rect 15059 5412 15115 5414
rect 15139 5412 15195 5414
rect 15219 5412 15275 5414
rect 14979 4378 15035 4380
rect 15059 4378 15115 4380
rect 15139 4378 15195 4380
rect 15219 4378 15275 4380
rect 14979 4326 15025 4378
rect 15025 4326 15035 4378
rect 15059 4326 15089 4378
rect 15089 4326 15101 4378
rect 15101 4326 15115 4378
rect 15139 4326 15153 4378
rect 15153 4326 15165 4378
rect 15165 4326 15195 4378
rect 15219 4326 15229 4378
rect 15229 4326 15275 4378
rect 14979 4324 15035 4326
rect 15059 4324 15115 4326
rect 15139 4324 15195 4326
rect 15219 4324 15275 4326
rect 10501 3834 10557 3836
rect 10581 3834 10637 3836
rect 10661 3834 10717 3836
rect 10741 3834 10797 3836
rect 10501 3782 10547 3834
rect 10547 3782 10557 3834
rect 10581 3782 10611 3834
rect 10611 3782 10623 3834
rect 10623 3782 10637 3834
rect 10661 3782 10675 3834
rect 10675 3782 10687 3834
rect 10687 3782 10717 3834
rect 10741 3782 10751 3834
rect 10751 3782 10797 3834
rect 10501 3780 10557 3782
rect 10581 3780 10637 3782
rect 10661 3780 10717 3782
rect 10741 3780 10797 3782
rect 14319 3834 14375 3836
rect 14399 3834 14455 3836
rect 14479 3834 14535 3836
rect 14559 3834 14615 3836
rect 14319 3782 14365 3834
rect 14365 3782 14375 3834
rect 14399 3782 14429 3834
rect 14429 3782 14441 3834
rect 14441 3782 14455 3834
rect 14479 3782 14493 3834
rect 14493 3782 14505 3834
rect 14505 3782 14535 3834
rect 14559 3782 14569 3834
rect 14569 3782 14615 3834
rect 14319 3780 14375 3782
rect 14399 3780 14455 3782
rect 14479 3780 14535 3782
rect 14559 3780 14615 3782
rect 15934 3440 15990 3496
rect 11161 3290 11217 3292
rect 11241 3290 11297 3292
rect 11321 3290 11377 3292
rect 11401 3290 11457 3292
rect 11161 3238 11207 3290
rect 11207 3238 11217 3290
rect 11241 3238 11271 3290
rect 11271 3238 11283 3290
rect 11283 3238 11297 3290
rect 11321 3238 11335 3290
rect 11335 3238 11347 3290
rect 11347 3238 11377 3290
rect 11401 3238 11411 3290
rect 11411 3238 11457 3290
rect 11161 3236 11217 3238
rect 11241 3236 11297 3238
rect 11321 3236 11377 3238
rect 11401 3236 11457 3238
rect 10501 2746 10557 2748
rect 10581 2746 10637 2748
rect 10661 2746 10717 2748
rect 10741 2746 10797 2748
rect 10501 2694 10547 2746
rect 10547 2694 10557 2746
rect 10581 2694 10611 2746
rect 10611 2694 10623 2746
rect 10623 2694 10637 2746
rect 10661 2694 10675 2746
rect 10675 2694 10687 2746
rect 10687 2694 10717 2746
rect 10741 2694 10751 2746
rect 10751 2694 10797 2746
rect 10501 2692 10557 2694
rect 10581 2692 10637 2694
rect 10661 2692 10717 2694
rect 10741 2692 10797 2694
rect 14979 3290 15035 3292
rect 15059 3290 15115 3292
rect 15139 3290 15195 3292
rect 15219 3290 15275 3292
rect 14979 3238 15025 3290
rect 15025 3238 15035 3290
rect 15059 3238 15089 3290
rect 15089 3238 15101 3290
rect 15101 3238 15115 3290
rect 15139 3238 15153 3290
rect 15153 3238 15165 3290
rect 15165 3238 15195 3290
rect 15219 3238 15229 3290
rect 15229 3238 15275 3290
rect 14979 3236 15035 3238
rect 15059 3236 15115 3238
rect 15139 3236 15195 3238
rect 15219 3236 15275 3238
rect 14319 2746 14375 2748
rect 14399 2746 14455 2748
rect 14479 2746 14535 2748
rect 14559 2746 14615 2748
rect 14319 2694 14365 2746
rect 14365 2694 14375 2746
rect 14399 2694 14429 2746
rect 14429 2694 14441 2746
rect 14441 2694 14455 2746
rect 14479 2694 14493 2746
rect 14493 2694 14505 2746
rect 14505 2694 14535 2746
rect 14559 2694 14569 2746
rect 14569 2694 14615 2746
rect 14319 2692 14375 2694
rect 14399 2692 14455 2694
rect 14479 2692 14535 2694
rect 14559 2692 14615 2694
rect 3525 2202 3581 2204
rect 3605 2202 3661 2204
rect 3685 2202 3741 2204
rect 3765 2202 3821 2204
rect 3525 2150 3571 2202
rect 3571 2150 3581 2202
rect 3605 2150 3635 2202
rect 3635 2150 3647 2202
rect 3647 2150 3661 2202
rect 3685 2150 3699 2202
rect 3699 2150 3711 2202
rect 3711 2150 3741 2202
rect 3765 2150 3775 2202
rect 3775 2150 3821 2202
rect 3525 2148 3581 2150
rect 3605 2148 3661 2150
rect 3685 2148 3741 2150
rect 3765 2148 3821 2150
rect 7343 2202 7399 2204
rect 7423 2202 7479 2204
rect 7503 2202 7559 2204
rect 7583 2202 7639 2204
rect 7343 2150 7389 2202
rect 7389 2150 7399 2202
rect 7423 2150 7453 2202
rect 7453 2150 7465 2202
rect 7465 2150 7479 2202
rect 7503 2150 7517 2202
rect 7517 2150 7529 2202
rect 7529 2150 7559 2202
rect 7583 2150 7593 2202
rect 7593 2150 7639 2202
rect 7343 2148 7399 2150
rect 7423 2148 7479 2150
rect 7503 2148 7559 2150
rect 7583 2148 7639 2150
rect 11161 2202 11217 2204
rect 11241 2202 11297 2204
rect 11321 2202 11377 2204
rect 11401 2202 11457 2204
rect 11161 2150 11207 2202
rect 11207 2150 11217 2202
rect 11241 2150 11271 2202
rect 11271 2150 11283 2202
rect 11283 2150 11297 2202
rect 11321 2150 11335 2202
rect 11335 2150 11347 2202
rect 11347 2150 11377 2202
rect 11401 2150 11411 2202
rect 11411 2150 11457 2202
rect 11161 2148 11217 2150
rect 11241 2148 11297 2150
rect 11321 2148 11377 2150
rect 11401 2148 11457 2150
rect 14979 2202 15035 2204
rect 15059 2202 15115 2204
rect 15139 2202 15195 2204
rect 15219 2202 15275 2204
rect 14979 2150 15025 2202
rect 15025 2150 15035 2202
rect 15059 2150 15089 2202
rect 15089 2150 15101 2202
rect 15101 2150 15115 2202
rect 15139 2150 15153 2202
rect 15153 2150 15165 2202
rect 15165 2150 15195 2202
rect 15219 2150 15229 2202
rect 15229 2150 15275 2202
rect 14979 2148 15035 2150
rect 15059 2148 15115 2150
rect 15139 2148 15195 2150
rect 15219 2148 15275 2150
<< metal3 >>
rect 3515 17440 3831 17441
rect 3515 17376 3521 17440
rect 3585 17376 3601 17440
rect 3665 17376 3681 17440
rect 3745 17376 3761 17440
rect 3825 17376 3831 17440
rect 3515 17375 3831 17376
rect 7333 17440 7649 17441
rect 7333 17376 7339 17440
rect 7403 17376 7419 17440
rect 7483 17376 7499 17440
rect 7563 17376 7579 17440
rect 7643 17376 7649 17440
rect 7333 17375 7649 17376
rect 11151 17440 11467 17441
rect 11151 17376 11157 17440
rect 11221 17376 11237 17440
rect 11301 17376 11317 17440
rect 11381 17376 11397 17440
rect 11461 17376 11467 17440
rect 11151 17375 11467 17376
rect 14969 17440 15285 17441
rect 14969 17376 14975 17440
rect 15039 17376 15055 17440
rect 15119 17376 15135 17440
rect 15199 17376 15215 17440
rect 15279 17376 15285 17440
rect 14969 17375 15285 17376
rect 2855 16896 3171 16897
rect 2855 16832 2861 16896
rect 2925 16832 2941 16896
rect 3005 16832 3021 16896
rect 3085 16832 3101 16896
rect 3165 16832 3171 16896
rect 2855 16831 3171 16832
rect 6673 16896 6989 16897
rect 6673 16832 6679 16896
rect 6743 16832 6759 16896
rect 6823 16832 6839 16896
rect 6903 16832 6919 16896
rect 6983 16832 6989 16896
rect 6673 16831 6989 16832
rect 10491 16896 10807 16897
rect 10491 16832 10497 16896
rect 10561 16832 10577 16896
rect 10641 16832 10657 16896
rect 10721 16832 10737 16896
rect 10801 16832 10807 16896
rect 10491 16831 10807 16832
rect 14309 16896 14625 16897
rect 14309 16832 14315 16896
rect 14379 16832 14395 16896
rect 14459 16832 14475 16896
rect 14539 16832 14555 16896
rect 14619 16832 14625 16896
rect 14309 16831 14625 16832
rect 3515 16352 3831 16353
rect 3515 16288 3521 16352
rect 3585 16288 3601 16352
rect 3665 16288 3681 16352
rect 3745 16288 3761 16352
rect 3825 16288 3831 16352
rect 3515 16287 3831 16288
rect 7333 16352 7649 16353
rect 7333 16288 7339 16352
rect 7403 16288 7419 16352
rect 7483 16288 7499 16352
rect 7563 16288 7579 16352
rect 7643 16288 7649 16352
rect 7333 16287 7649 16288
rect 11151 16352 11467 16353
rect 11151 16288 11157 16352
rect 11221 16288 11237 16352
rect 11301 16288 11317 16352
rect 11381 16288 11397 16352
rect 11461 16288 11467 16352
rect 11151 16287 11467 16288
rect 14969 16352 15285 16353
rect 14969 16288 14975 16352
rect 15039 16288 15055 16352
rect 15119 16288 15135 16352
rect 15199 16288 15215 16352
rect 15279 16288 15285 16352
rect 14969 16287 15285 16288
rect 2855 15808 3171 15809
rect 2855 15744 2861 15808
rect 2925 15744 2941 15808
rect 3005 15744 3021 15808
rect 3085 15744 3101 15808
rect 3165 15744 3171 15808
rect 2855 15743 3171 15744
rect 6673 15808 6989 15809
rect 6673 15744 6679 15808
rect 6743 15744 6759 15808
rect 6823 15744 6839 15808
rect 6903 15744 6919 15808
rect 6983 15744 6989 15808
rect 6673 15743 6989 15744
rect 10491 15808 10807 15809
rect 10491 15744 10497 15808
rect 10561 15744 10577 15808
rect 10641 15744 10657 15808
rect 10721 15744 10737 15808
rect 10801 15744 10807 15808
rect 10491 15743 10807 15744
rect 14309 15808 14625 15809
rect 14309 15744 14315 15808
rect 14379 15744 14395 15808
rect 14459 15744 14475 15808
rect 14539 15744 14555 15808
rect 14619 15744 14625 15808
rect 14309 15743 14625 15744
rect 3515 15264 3831 15265
rect 3515 15200 3521 15264
rect 3585 15200 3601 15264
rect 3665 15200 3681 15264
rect 3745 15200 3761 15264
rect 3825 15200 3831 15264
rect 3515 15199 3831 15200
rect 7333 15264 7649 15265
rect 7333 15200 7339 15264
rect 7403 15200 7419 15264
rect 7483 15200 7499 15264
rect 7563 15200 7579 15264
rect 7643 15200 7649 15264
rect 7333 15199 7649 15200
rect 11151 15264 11467 15265
rect 11151 15200 11157 15264
rect 11221 15200 11237 15264
rect 11301 15200 11317 15264
rect 11381 15200 11397 15264
rect 11461 15200 11467 15264
rect 11151 15199 11467 15200
rect 14969 15264 15285 15265
rect 14969 15200 14975 15264
rect 15039 15200 15055 15264
rect 15119 15200 15135 15264
rect 15199 15200 15215 15264
rect 15279 15200 15285 15264
rect 14969 15199 15285 15200
rect 16021 15058 16087 15061
rect 16699 15058 17499 15088
rect 16021 15056 17499 15058
rect 16021 15000 16026 15056
rect 16082 15000 17499 15056
rect 16021 14998 17499 15000
rect 16021 14995 16087 14998
rect 16699 14968 17499 14998
rect 2855 14720 3171 14721
rect 2855 14656 2861 14720
rect 2925 14656 2941 14720
rect 3005 14656 3021 14720
rect 3085 14656 3101 14720
rect 3165 14656 3171 14720
rect 2855 14655 3171 14656
rect 6673 14720 6989 14721
rect 6673 14656 6679 14720
rect 6743 14656 6759 14720
rect 6823 14656 6839 14720
rect 6903 14656 6919 14720
rect 6983 14656 6989 14720
rect 6673 14655 6989 14656
rect 10491 14720 10807 14721
rect 10491 14656 10497 14720
rect 10561 14656 10577 14720
rect 10641 14656 10657 14720
rect 10721 14656 10737 14720
rect 10801 14656 10807 14720
rect 10491 14655 10807 14656
rect 14309 14720 14625 14721
rect 14309 14656 14315 14720
rect 14379 14656 14395 14720
rect 14459 14656 14475 14720
rect 14539 14656 14555 14720
rect 14619 14656 14625 14720
rect 14309 14655 14625 14656
rect 0 14378 800 14408
rect 933 14378 999 14381
rect 0 14376 999 14378
rect 0 14320 938 14376
rect 994 14320 999 14376
rect 0 14318 999 14320
rect 0 14288 800 14318
rect 933 14315 999 14318
rect 3515 14176 3831 14177
rect 3515 14112 3521 14176
rect 3585 14112 3601 14176
rect 3665 14112 3681 14176
rect 3745 14112 3761 14176
rect 3825 14112 3831 14176
rect 3515 14111 3831 14112
rect 7333 14176 7649 14177
rect 7333 14112 7339 14176
rect 7403 14112 7419 14176
rect 7483 14112 7499 14176
rect 7563 14112 7579 14176
rect 7643 14112 7649 14176
rect 7333 14111 7649 14112
rect 11151 14176 11467 14177
rect 11151 14112 11157 14176
rect 11221 14112 11237 14176
rect 11301 14112 11317 14176
rect 11381 14112 11397 14176
rect 11461 14112 11467 14176
rect 11151 14111 11467 14112
rect 14969 14176 15285 14177
rect 14969 14112 14975 14176
rect 15039 14112 15055 14176
rect 15119 14112 15135 14176
rect 15199 14112 15215 14176
rect 15279 14112 15285 14176
rect 14969 14111 15285 14112
rect 2855 13632 3171 13633
rect 2855 13568 2861 13632
rect 2925 13568 2941 13632
rect 3005 13568 3021 13632
rect 3085 13568 3101 13632
rect 3165 13568 3171 13632
rect 2855 13567 3171 13568
rect 6673 13632 6989 13633
rect 6673 13568 6679 13632
rect 6743 13568 6759 13632
rect 6823 13568 6839 13632
rect 6903 13568 6919 13632
rect 6983 13568 6989 13632
rect 6673 13567 6989 13568
rect 10491 13632 10807 13633
rect 10491 13568 10497 13632
rect 10561 13568 10577 13632
rect 10641 13568 10657 13632
rect 10721 13568 10737 13632
rect 10801 13568 10807 13632
rect 10491 13567 10807 13568
rect 14309 13632 14625 13633
rect 14309 13568 14315 13632
rect 14379 13568 14395 13632
rect 14459 13568 14475 13632
rect 14539 13568 14555 13632
rect 14619 13568 14625 13632
rect 14309 13567 14625 13568
rect 3515 13088 3831 13089
rect 0 13018 800 13048
rect 3515 13024 3521 13088
rect 3585 13024 3601 13088
rect 3665 13024 3681 13088
rect 3745 13024 3761 13088
rect 3825 13024 3831 13088
rect 3515 13023 3831 13024
rect 7333 13088 7649 13089
rect 7333 13024 7339 13088
rect 7403 13024 7419 13088
rect 7483 13024 7499 13088
rect 7563 13024 7579 13088
rect 7643 13024 7649 13088
rect 7333 13023 7649 13024
rect 11151 13088 11467 13089
rect 11151 13024 11157 13088
rect 11221 13024 11237 13088
rect 11301 13024 11317 13088
rect 11381 13024 11397 13088
rect 11461 13024 11467 13088
rect 11151 13023 11467 13024
rect 14969 13088 15285 13089
rect 14969 13024 14975 13088
rect 15039 13024 15055 13088
rect 15119 13024 15135 13088
rect 15199 13024 15215 13088
rect 15279 13024 15285 13088
rect 14969 13023 15285 13024
rect 933 13018 999 13021
rect 0 13016 999 13018
rect 0 12960 938 13016
rect 994 12960 999 13016
rect 0 12958 999 12960
rect 0 12928 800 12958
rect 933 12955 999 12958
rect 15929 13018 15995 13021
rect 16699 13018 17499 13048
rect 15929 13016 17499 13018
rect 15929 12960 15934 13016
rect 15990 12960 17499 13016
rect 15929 12958 17499 12960
rect 15929 12955 15995 12958
rect 16699 12928 17499 12958
rect 2855 12544 3171 12545
rect 2855 12480 2861 12544
rect 2925 12480 2941 12544
rect 3005 12480 3021 12544
rect 3085 12480 3101 12544
rect 3165 12480 3171 12544
rect 2855 12479 3171 12480
rect 6673 12544 6989 12545
rect 6673 12480 6679 12544
rect 6743 12480 6759 12544
rect 6823 12480 6839 12544
rect 6903 12480 6919 12544
rect 6983 12480 6989 12544
rect 6673 12479 6989 12480
rect 10491 12544 10807 12545
rect 10491 12480 10497 12544
rect 10561 12480 10577 12544
rect 10641 12480 10657 12544
rect 10721 12480 10737 12544
rect 10801 12480 10807 12544
rect 10491 12479 10807 12480
rect 14309 12544 14625 12545
rect 14309 12480 14315 12544
rect 14379 12480 14395 12544
rect 14459 12480 14475 12544
rect 14539 12480 14555 12544
rect 14619 12480 14625 12544
rect 14309 12479 14625 12480
rect 0 12338 800 12368
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12248 800 12278
rect 1393 12275 1459 12278
rect 3515 12000 3831 12001
rect 3515 11936 3521 12000
rect 3585 11936 3601 12000
rect 3665 11936 3681 12000
rect 3745 11936 3761 12000
rect 3825 11936 3831 12000
rect 3515 11935 3831 11936
rect 7333 12000 7649 12001
rect 7333 11936 7339 12000
rect 7403 11936 7419 12000
rect 7483 11936 7499 12000
rect 7563 11936 7579 12000
rect 7643 11936 7649 12000
rect 7333 11935 7649 11936
rect 11151 12000 11467 12001
rect 11151 11936 11157 12000
rect 11221 11936 11237 12000
rect 11301 11936 11317 12000
rect 11381 11936 11397 12000
rect 11461 11936 11467 12000
rect 11151 11935 11467 11936
rect 14969 12000 15285 12001
rect 14969 11936 14975 12000
rect 15039 11936 15055 12000
rect 15119 11936 15135 12000
rect 15199 11936 15215 12000
rect 15279 11936 15285 12000
rect 14969 11935 15285 11936
rect 2855 11456 3171 11457
rect 2855 11392 2861 11456
rect 2925 11392 2941 11456
rect 3005 11392 3021 11456
rect 3085 11392 3101 11456
rect 3165 11392 3171 11456
rect 2855 11391 3171 11392
rect 6673 11456 6989 11457
rect 6673 11392 6679 11456
rect 6743 11392 6759 11456
rect 6823 11392 6839 11456
rect 6903 11392 6919 11456
rect 6983 11392 6989 11456
rect 6673 11391 6989 11392
rect 10491 11456 10807 11457
rect 10491 11392 10497 11456
rect 10561 11392 10577 11456
rect 10641 11392 10657 11456
rect 10721 11392 10737 11456
rect 10801 11392 10807 11456
rect 10491 11391 10807 11392
rect 14309 11456 14625 11457
rect 14309 11392 14315 11456
rect 14379 11392 14395 11456
rect 14459 11392 14475 11456
rect 14539 11392 14555 11456
rect 14619 11392 14625 11456
rect 14309 11391 14625 11392
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 16021 10978 16087 10981
rect 16699 10978 17499 11008
rect 16021 10976 17499 10978
rect 16021 10920 16026 10976
rect 16082 10920 17499 10976
rect 16021 10918 17499 10920
rect 16021 10915 16087 10918
rect 3515 10912 3831 10913
rect 3515 10848 3521 10912
rect 3585 10848 3601 10912
rect 3665 10848 3681 10912
rect 3745 10848 3761 10912
rect 3825 10848 3831 10912
rect 3515 10847 3831 10848
rect 7333 10912 7649 10913
rect 7333 10848 7339 10912
rect 7403 10848 7419 10912
rect 7483 10848 7499 10912
rect 7563 10848 7579 10912
rect 7643 10848 7649 10912
rect 7333 10847 7649 10848
rect 11151 10912 11467 10913
rect 11151 10848 11157 10912
rect 11221 10848 11237 10912
rect 11301 10848 11317 10912
rect 11381 10848 11397 10912
rect 11461 10848 11467 10912
rect 11151 10847 11467 10848
rect 14969 10912 15285 10913
rect 14969 10848 14975 10912
rect 15039 10848 15055 10912
rect 15119 10848 15135 10912
rect 15199 10848 15215 10912
rect 15279 10848 15285 10912
rect 16699 10888 17499 10918
rect 14969 10847 15285 10848
rect 2855 10368 3171 10369
rect 0 10298 800 10328
rect 2855 10304 2861 10368
rect 2925 10304 2941 10368
rect 3005 10304 3021 10368
rect 3085 10304 3101 10368
rect 3165 10304 3171 10368
rect 2855 10303 3171 10304
rect 6673 10368 6989 10369
rect 6673 10304 6679 10368
rect 6743 10304 6759 10368
rect 6823 10304 6839 10368
rect 6903 10304 6919 10368
rect 6983 10304 6989 10368
rect 6673 10303 6989 10304
rect 10491 10368 10807 10369
rect 10491 10304 10497 10368
rect 10561 10304 10577 10368
rect 10641 10304 10657 10368
rect 10721 10304 10737 10368
rect 10801 10304 10807 10368
rect 10491 10303 10807 10304
rect 14309 10368 14625 10369
rect 14309 10304 14315 10368
rect 14379 10304 14395 10368
rect 14459 10304 14475 10368
rect 14539 10304 14555 10368
rect 14619 10304 14625 10368
rect 14309 10303 14625 10304
rect 933 10298 999 10301
rect 0 10296 999 10298
rect 0 10240 938 10296
rect 994 10240 999 10296
rect 0 10238 999 10240
rect 0 10208 800 10238
rect 933 10235 999 10238
rect 3515 9824 3831 9825
rect 3515 9760 3521 9824
rect 3585 9760 3601 9824
rect 3665 9760 3681 9824
rect 3745 9760 3761 9824
rect 3825 9760 3831 9824
rect 3515 9759 3831 9760
rect 7333 9824 7649 9825
rect 7333 9760 7339 9824
rect 7403 9760 7419 9824
rect 7483 9760 7499 9824
rect 7563 9760 7579 9824
rect 7643 9760 7649 9824
rect 7333 9759 7649 9760
rect 11151 9824 11467 9825
rect 11151 9760 11157 9824
rect 11221 9760 11237 9824
rect 11301 9760 11317 9824
rect 11381 9760 11397 9824
rect 11461 9760 11467 9824
rect 11151 9759 11467 9760
rect 14969 9824 15285 9825
rect 14969 9760 14975 9824
rect 15039 9760 15055 9824
rect 15119 9760 15135 9824
rect 15199 9760 15215 9824
rect 15279 9760 15285 9824
rect 14969 9759 15285 9760
rect 0 9618 800 9648
rect 1485 9618 1551 9621
rect 0 9616 1551 9618
rect 0 9560 1490 9616
rect 1546 9560 1551 9616
rect 0 9558 1551 9560
rect 0 9528 800 9558
rect 1485 9555 1551 9558
rect 7465 9618 7531 9621
rect 9029 9618 9095 9621
rect 7465 9616 9095 9618
rect 7465 9560 7470 9616
rect 7526 9560 9034 9616
rect 9090 9560 9095 9616
rect 7465 9558 9095 9560
rect 7465 9555 7531 9558
rect 9029 9555 9095 9558
rect 16021 9618 16087 9621
rect 16699 9618 17499 9648
rect 16021 9616 17499 9618
rect 16021 9560 16026 9616
rect 16082 9560 17499 9616
rect 16021 9558 17499 9560
rect 16021 9555 16087 9558
rect 16699 9528 17499 9558
rect 2855 9280 3171 9281
rect 2855 9216 2861 9280
rect 2925 9216 2941 9280
rect 3005 9216 3021 9280
rect 3085 9216 3101 9280
rect 3165 9216 3171 9280
rect 2855 9215 3171 9216
rect 6673 9280 6989 9281
rect 6673 9216 6679 9280
rect 6743 9216 6759 9280
rect 6823 9216 6839 9280
rect 6903 9216 6919 9280
rect 6983 9216 6989 9280
rect 6673 9215 6989 9216
rect 10491 9280 10807 9281
rect 10491 9216 10497 9280
rect 10561 9216 10577 9280
rect 10641 9216 10657 9280
rect 10721 9216 10737 9280
rect 10801 9216 10807 9280
rect 10491 9215 10807 9216
rect 14309 9280 14625 9281
rect 14309 9216 14315 9280
rect 14379 9216 14395 9280
rect 14459 9216 14475 9280
rect 14539 9216 14555 9280
rect 14619 9216 14625 9280
rect 14309 9215 14625 9216
rect 7465 9074 7531 9077
rect 8385 9074 8451 9077
rect 7465 9072 8451 9074
rect 7465 9016 7470 9072
rect 7526 9016 8390 9072
rect 8446 9016 8451 9072
rect 7465 9014 8451 9016
rect 7465 9011 7531 9014
rect 8385 9011 8451 9014
rect 0 8938 800 8968
rect 933 8938 999 8941
rect 0 8936 999 8938
rect 0 8880 938 8936
rect 994 8880 999 8936
rect 0 8878 999 8880
rect 0 8848 800 8878
rect 933 8875 999 8878
rect 3515 8736 3831 8737
rect 3515 8672 3521 8736
rect 3585 8672 3601 8736
rect 3665 8672 3681 8736
rect 3745 8672 3761 8736
rect 3825 8672 3831 8736
rect 3515 8671 3831 8672
rect 7333 8736 7649 8737
rect 7333 8672 7339 8736
rect 7403 8672 7419 8736
rect 7483 8672 7499 8736
rect 7563 8672 7579 8736
rect 7643 8672 7649 8736
rect 7333 8671 7649 8672
rect 11151 8736 11467 8737
rect 11151 8672 11157 8736
rect 11221 8672 11237 8736
rect 11301 8672 11317 8736
rect 11381 8672 11397 8736
rect 11461 8672 11467 8736
rect 11151 8671 11467 8672
rect 14969 8736 15285 8737
rect 14969 8672 14975 8736
rect 15039 8672 15055 8736
rect 15119 8672 15135 8736
rect 15199 8672 15215 8736
rect 15279 8672 15285 8736
rect 14969 8671 15285 8672
rect 0 8258 800 8288
rect 2681 8258 2747 8261
rect 0 8256 2747 8258
rect 0 8200 2686 8256
rect 2742 8200 2747 8256
rect 0 8198 2747 8200
rect 0 8168 800 8198
rect 2681 8195 2747 8198
rect 2855 8192 3171 8193
rect 2855 8128 2861 8192
rect 2925 8128 2941 8192
rect 3005 8128 3021 8192
rect 3085 8128 3101 8192
rect 3165 8128 3171 8192
rect 2855 8127 3171 8128
rect 6673 8192 6989 8193
rect 6673 8128 6679 8192
rect 6743 8128 6759 8192
rect 6823 8128 6839 8192
rect 6903 8128 6919 8192
rect 6983 8128 6989 8192
rect 6673 8127 6989 8128
rect 10491 8192 10807 8193
rect 10491 8128 10497 8192
rect 10561 8128 10577 8192
rect 10641 8128 10657 8192
rect 10721 8128 10737 8192
rect 10801 8128 10807 8192
rect 10491 8127 10807 8128
rect 14309 8192 14625 8193
rect 14309 8128 14315 8192
rect 14379 8128 14395 8192
rect 14459 8128 14475 8192
rect 14539 8128 14555 8192
rect 14619 8128 14625 8192
rect 14309 8127 14625 8128
rect 2497 7850 2563 7853
rect 4337 7850 4403 7853
rect 2497 7848 4403 7850
rect 2497 7792 2502 7848
rect 2558 7792 4342 7848
rect 4398 7792 4403 7848
rect 2497 7790 4403 7792
rect 2497 7787 2563 7790
rect 4337 7787 4403 7790
rect 3515 7648 3831 7649
rect 0 7578 800 7608
rect 3515 7584 3521 7648
rect 3585 7584 3601 7648
rect 3665 7584 3681 7648
rect 3745 7584 3761 7648
rect 3825 7584 3831 7648
rect 3515 7583 3831 7584
rect 7333 7648 7649 7649
rect 7333 7584 7339 7648
rect 7403 7584 7419 7648
rect 7483 7584 7499 7648
rect 7563 7584 7579 7648
rect 7643 7584 7649 7648
rect 7333 7583 7649 7584
rect 11151 7648 11467 7649
rect 11151 7584 11157 7648
rect 11221 7584 11237 7648
rect 11301 7584 11317 7648
rect 11381 7584 11397 7648
rect 11461 7584 11467 7648
rect 11151 7583 11467 7584
rect 14969 7648 15285 7649
rect 14969 7584 14975 7648
rect 15039 7584 15055 7648
rect 15119 7584 15135 7648
rect 15199 7584 15215 7648
rect 15279 7584 15285 7648
rect 14969 7583 15285 7584
rect 933 7578 999 7581
rect 0 7576 999 7578
rect 0 7520 938 7576
rect 994 7520 999 7576
rect 0 7518 999 7520
rect 0 7488 800 7518
rect 933 7515 999 7518
rect 15929 7578 15995 7581
rect 16699 7578 17499 7608
rect 15929 7576 17499 7578
rect 15929 7520 15934 7576
rect 15990 7520 17499 7576
rect 15929 7518 17499 7520
rect 15929 7515 15995 7518
rect 16699 7488 17499 7518
rect 4245 7306 4311 7309
rect 5441 7306 5507 7309
rect 4245 7304 5507 7306
rect 4245 7248 4250 7304
rect 4306 7248 5446 7304
rect 5502 7248 5507 7304
rect 4245 7246 5507 7248
rect 4245 7243 4311 7246
rect 5441 7243 5507 7246
rect 2855 7104 3171 7105
rect 2855 7040 2861 7104
rect 2925 7040 2941 7104
rect 3005 7040 3021 7104
rect 3085 7040 3101 7104
rect 3165 7040 3171 7104
rect 2855 7039 3171 7040
rect 6673 7104 6989 7105
rect 6673 7040 6679 7104
rect 6743 7040 6759 7104
rect 6823 7040 6839 7104
rect 6903 7040 6919 7104
rect 6983 7040 6989 7104
rect 6673 7039 6989 7040
rect 10491 7104 10807 7105
rect 10491 7040 10497 7104
rect 10561 7040 10577 7104
rect 10641 7040 10657 7104
rect 10721 7040 10737 7104
rect 10801 7040 10807 7104
rect 10491 7039 10807 7040
rect 14309 7104 14625 7105
rect 14309 7040 14315 7104
rect 14379 7040 14395 7104
rect 14459 7040 14475 7104
rect 14539 7040 14555 7104
rect 14619 7040 14625 7104
rect 14309 7039 14625 7040
rect 0 6898 800 6928
rect 933 6898 999 6901
rect 0 6896 999 6898
rect 0 6840 938 6896
rect 994 6840 999 6896
rect 0 6838 999 6840
rect 0 6808 800 6838
rect 933 6835 999 6838
rect 3515 6560 3831 6561
rect 3515 6496 3521 6560
rect 3585 6496 3601 6560
rect 3665 6496 3681 6560
rect 3745 6496 3761 6560
rect 3825 6496 3831 6560
rect 3515 6495 3831 6496
rect 7333 6560 7649 6561
rect 7333 6496 7339 6560
rect 7403 6496 7419 6560
rect 7483 6496 7499 6560
rect 7563 6496 7579 6560
rect 7643 6496 7649 6560
rect 7333 6495 7649 6496
rect 11151 6560 11467 6561
rect 11151 6496 11157 6560
rect 11221 6496 11237 6560
rect 11301 6496 11317 6560
rect 11381 6496 11397 6560
rect 11461 6496 11467 6560
rect 11151 6495 11467 6496
rect 14969 6560 15285 6561
rect 14969 6496 14975 6560
rect 15039 6496 15055 6560
rect 15119 6496 15135 6560
rect 15199 6496 15215 6560
rect 15279 6496 15285 6560
rect 14969 6495 15285 6496
rect 0 6218 800 6248
rect 2773 6218 2839 6221
rect 0 6216 2839 6218
rect 0 6160 2778 6216
rect 2834 6160 2839 6216
rect 0 6158 2839 6160
rect 0 6128 800 6158
rect 2773 6155 2839 6158
rect 2855 6016 3171 6017
rect 2855 5952 2861 6016
rect 2925 5952 2941 6016
rect 3005 5952 3021 6016
rect 3085 5952 3101 6016
rect 3165 5952 3171 6016
rect 2855 5951 3171 5952
rect 6673 6016 6989 6017
rect 6673 5952 6679 6016
rect 6743 5952 6759 6016
rect 6823 5952 6839 6016
rect 6903 5952 6919 6016
rect 6983 5952 6989 6016
rect 6673 5951 6989 5952
rect 10491 6016 10807 6017
rect 10491 5952 10497 6016
rect 10561 5952 10577 6016
rect 10641 5952 10657 6016
rect 10721 5952 10737 6016
rect 10801 5952 10807 6016
rect 10491 5951 10807 5952
rect 14309 6016 14625 6017
rect 14309 5952 14315 6016
rect 14379 5952 14395 6016
rect 14459 5952 14475 6016
rect 14539 5952 14555 6016
rect 14619 5952 14625 6016
rect 14309 5951 14625 5952
rect 0 5538 800 5568
rect 933 5538 999 5541
rect 0 5536 999 5538
rect 0 5480 938 5536
rect 994 5480 999 5536
rect 0 5478 999 5480
rect 0 5448 800 5478
rect 933 5475 999 5478
rect 16021 5538 16087 5541
rect 16699 5538 17499 5568
rect 16021 5536 17499 5538
rect 16021 5480 16026 5536
rect 16082 5480 17499 5536
rect 16021 5478 17499 5480
rect 16021 5475 16087 5478
rect 3515 5472 3831 5473
rect 3515 5408 3521 5472
rect 3585 5408 3601 5472
rect 3665 5408 3681 5472
rect 3745 5408 3761 5472
rect 3825 5408 3831 5472
rect 3515 5407 3831 5408
rect 7333 5472 7649 5473
rect 7333 5408 7339 5472
rect 7403 5408 7419 5472
rect 7483 5408 7499 5472
rect 7563 5408 7579 5472
rect 7643 5408 7649 5472
rect 7333 5407 7649 5408
rect 11151 5472 11467 5473
rect 11151 5408 11157 5472
rect 11221 5408 11237 5472
rect 11301 5408 11317 5472
rect 11381 5408 11397 5472
rect 11461 5408 11467 5472
rect 11151 5407 11467 5408
rect 14969 5472 15285 5473
rect 14969 5408 14975 5472
rect 15039 5408 15055 5472
rect 15119 5408 15135 5472
rect 15199 5408 15215 5472
rect 15279 5408 15285 5472
rect 16699 5448 17499 5478
rect 14969 5407 15285 5408
rect 2855 4928 3171 4929
rect 0 4858 800 4888
rect 2855 4864 2861 4928
rect 2925 4864 2941 4928
rect 3005 4864 3021 4928
rect 3085 4864 3101 4928
rect 3165 4864 3171 4928
rect 2855 4863 3171 4864
rect 6673 4928 6989 4929
rect 6673 4864 6679 4928
rect 6743 4864 6759 4928
rect 6823 4864 6839 4928
rect 6903 4864 6919 4928
rect 6983 4864 6989 4928
rect 6673 4863 6989 4864
rect 10491 4928 10807 4929
rect 10491 4864 10497 4928
rect 10561 4864 10577 4928
rect 10641 4864 10657 4928
rect 10721 4864 10737 4928
rect 10801 4864 10807 4928
rect 10491 4863 10807 4864
rect 14309 4928 14625 4929
rect 14309 4864 14315 4928
rect 14379 4864 14395 4928
rect 14459 4864 14475 4928
rect 14539 4864 14555 4928
rect 14619 4864 14625 4928
rect 14309 4863 14625 4864
rect 0 4798 1042 4858
rect 0 4768 800 4798
rect 982 4722 1042 4798
rect 1393 4722 1459 4725
rect 982 4720 1459 4722
rect 982 4664 1398 4720
rect 1454 4664 1459 4720
rect 982 4662 1459 4664
rect 1393 4659 1459 4662
rect 3515 4384 3831 4385
rect 3515 4320 3521 4384
rect 3585 4320 3601 4384
rect 3665 4320 3681 4384
rect 3745 4320 3761 4384
rect 3825 4320 3831 4384
rect 3515 4319 3831 4320
rect 7333 4384 7649 4385
rect 7333 4320 7339 4384
rect 7403 4320 7419 4384
rect 7483 4320 7499 4384
rect 7563 4320 7579 4384
rect 7643 4320 7649 4384
rect 7333 4319 7649 4320
rect 11151 4384 11467 4385
rect 11151 4320 11157 4384
rect 11221 4320 11237 4384
rect 11301 4320 11317 4384
rect 11381 4320 11397 4384
rect 11461 4320 11467 4384
rect 11151 4319 11467 4320
rect 14969 4384 15285 4385
rect 14969 4320 14975 4384
rect 15039 4320 15055 4384
rect 15119 4320 15135 4384
rect 15199 4320 15215 4384
rect 15279 4320 15285 4384
rect 14969 4319 15285 4320
rect 0 4178 800 4208
rect 1025 4178 1091 4181
rect 0 4176 1091 4178
rect 0 4120 1030 4176
rect 1086 4120 1091 4176
rect 0 4118 1091 4120
rect 0 4088 800 4118
rect 1025 4115 1091 4118
rect 2855 3840 3171 3841
rect 2855 3776 2861 3840
rect 2925 3776 2941 3840
rect 3005 3776 3021 3840
rect 3085 3776 3101 3840
rect 3165 3776 3171 3840
rect 2855 3775 3171 3776
rect 6673 3840 6989 3841
rect 6673 3776 6679 3840
rect 6743 3776 6759 3840
rect 6823 3776 6839 3840
rect 6903 3776 6919 3840
rect 6983 3776 6989 3840
rect 6673 3775 6989 3776
rect 10491 3840 10807 3841
rect 10491 3776 10497 3840
rect 10561 3776 10577 3840
rect 10641 3776 10657 3840
rect 10721 3776 10737 3840
rect 10801 3776 10807 3840
rect 10491 3775 10807 3776
rect 14309 3840 14625 3841
rect 14309 3776 14315 3840
rect 14379 3776 14395 3840
rect 14459 3776 14475 3840
rect 14539 3776 14555 3840
rect 14619 3776 14625 3840
rect 14309 3775 14625 3776
rect 6085 3634 6151 3637
rect 6729 3634 6795 3637
rect 6085 3632 6795 3634
rect 6085 3576 6090 3632
rect 6146 3576 6734 3632
rect 6790 3576 6795 3632
rect 6085 3574 6795 3576
rect 6085 3571 6151 3574
rect 6729 3571 6795 3574
rect 0 3498 800 3528
rect 933 3498 999 3501
rect 0 3496 999 3498
rect 0 3440 938 3496
rect 994 3440 999 3496
rect 0 3438 999 3440
rect 0 3408 800 3438
rect 933 3435 999 3438
rect 15929 3498 15995 3501
rect 16699 3498 17499 3528
rect 15929 3496 17499 3498
rect 15929 3440 15934 3496
rect 15990 3440 17499 3496
rect 15929 3438 17499 3440
rect 15929 3435 15995 3438
rect 16699 3408 17499 3438
rect 3515 3296 3831 3297
rect 3515 3232 3521 3296
rect 3585 3232 3601 3296
rect 3665 3232 3681 3296
rect 3745 3232 3761 3296
rect 3825 3232 3831 3296
rect 3515 3231 3831 3232
rect 7333 3296 7649 3297
rect 7333 3232 7339 3296
rect 7403 3232 7419 3296
rect 7483 3232 7499 3296
rect 7563 3232 7579 3296
rect 7643 3232 7649 3296
rect 7333 3231 7649 3232
rect 11151 3296 11467 3297
rect 11151 3232 11157 3296
rect 11221 3232 11237 3296
rect 11301 3232 11317 3296
rect 11381 3232 11397 3296
rect 11461 3232 11467 3296
rect 11151 3231 11467 3232
rect 14969 3296 15285 3297
rect 14969 3232 14975 3296
rect 15039 3232 15055 3296
rect 15119 3232 15135 3296
rect 15199 3232 15215 3296
rect 15279 3232 15285 3296
rect 14969 3231 15285 3232
rect 0 2818 800 2848
rect 933 2818 999 2821
rect 0 2816 999 2818
rect 0 2760 938 2816
rect 994 2760 999 2816
rect 0 2758 999 2760
rect 0 2728 800 2758
rect 933 2755 999 2758
rect 2855 2752 3171 2753
rect 2855 2688 2861 2752
rect 2925 2688 2941 2752
rect 3005 2688 3021 2752
rect 3085 2688 3101 2752
rect 3165 2688 3171 2752
rect 2855 2687 3171 2688
rect 6673 2752 6989 2753
rect 6673 2688 6679 2752
rect 6743 2688 6759 2752
rect 6823 2688 6839 2752
rect 6903 2688 6919 2752
rect 6983 2688 6989 2752
rect 6673 2687 6989 2688
rect 10491 2752 10807 2753
rect 10491 2688 10497 2752
rect 10561 2688 10577 2752
rect 10641 2688 10657 2752
rect 10721 2688 10737 2752
rect 10801 2688 10807 2752
rect 10491 2687 10807 2688
rect 14309 2752 14625 2753
rect 14309 2688 14315 2752
rect 14379 2688 14395 2752
rect 14459 2688 14475 2752
rect 14539 2688 14555 2752
rect 14619 2688 14625 2752
rect 14309 2687 14625 2688
rect 3515 2208 3831 2209
rect 3515 2144 3521 2208
rect 3585 2144 3601 2208
rect 3665 2144 3681 2208
rect 3745 2144 3761 2208
rect 3825 2144 3831 2208
rect 3515 2143 3831 2144
rect 7333 2208 7649 2209
rect 7333 2144 7339 2208
rect 7403 2144 7419 2208
rect 7483 2144 7499 2208
rect 7563 2144 7579 2208
rect 7643 2144 7649 2208
rect 7333 2143 7649 2144
rect 11151 2208 11467 2209
rect 11151 2144 11157 2208
rect 11221 2144 11237 2208
rect 11301 2144 11317 2208
rect 11381 2144 11397 2208
rect 11461 2144 11467 2208
rect 11151 2143 11467 2144
rect 14969 2208 15285 2209
rect 14969 2144 14975 2208
rect 15039 2144 15055 2208
rect 15119 2144 15135 2208
rect 15199 2144 15215 2208
rect 15279 2144 15285 2208
rect 14969 2143 15285 2144
<< via3 >>
rect 3521 17436 3585 17440
rect 3521 17380 3525 17436
rect 3525 17380 3581 17436
rect 3581 17380 3585 17436
rect 3521 17376 3585 17380
rect 3601 17436 3665 17440
rect 3601 17380 3605 17436
rect 3605 17380 3661 17436
rect 3661 17380 3665 17436
rect 3601 17376 3665 17380
rect 3681 17436 3745 17440
rect 3681 17380 3685 17436
rect 3685 17380 3741 17436
rect 3741 17380 3745 17436
rect 3681 17376 3745 17380
rect 3761 17436 3825 17440
rect 3761 17380 3765 17436
rect 3765 17380 3821 17436
rect 3821 17380 3825 17436
rect 3761 17376 3825 17380
rect 7339 17436 7403 17440
rect 7339 17380 7343 17436
rect 7343 17380 7399 17436
rect 7399 17380 7403 17436
rect 7339 17376 7403 17380
rect 7419 17436 7483 17440
rect 7419 17380 7423 17436
rect 7423 17380 7479 17436
rect 7479 17380 7483 17436
rect 7419 17376 7483 17380
rect 7499 17436 7563 17440
rect 7499 17380 7503 17436
rect 7503 17380 7559 17436
rect 7559 17380 7563 17436
rect 7499 17376 7563 17380
rect 7579 17436 7643 17440
rect 7579 17380 7583 17436
rect 7583 17380 7639 17436
rect 7639 17380 7643 17436
rect 7579 17376 7643 17380
rect 11157 17436 11221 17440
rect 11157 17380 11161 17436
rect 11161 17380 11217 17436
rect 11217 17380 11221 17436
rect 11157 17376 11221 17380
rect 11237 17436 11301 17440
rect 11237 17380 11241 17436
rect 11241 17380 11297 17436
rect 11297 17380 11301 17436
rect 11237 17376 11301 17380
rect 11317 17436 11381 17440
rect 11317 17380 11321 17436
rect 11321 17380 11377 17436
rect 11377 17380 11381 17436
rect 11317 17376 11381 17380
rect 11397 17436 11461 17440
rect 11397 17380 11401 17436
rect 11401 17380 11457 17436
rect 11457 17380 11461 17436
rect 11397 17376 11461 17380
rect 14975 17436 15039 17440
rect 14975 17380 14979 17436
rect 14979 17380 15035 17436
rect 15035 17380 15039 17436
rect 14975 17376 15039 17380
rect 15055 17436 15119 17440
rect 15055 17380 15059 17436
rect 15059 17380 15115 17436
rect 15115 17380 15119 17436
rect 15055 17376 15119 17380
rect 15135 17436 15199 17440
rect 15135 17380 15139 17436
rect 15139 17380 15195 17436
rect 15195 17380 15199 17436
rect 15135 17376 15199 17380
rect 15215 17436 15279 17440
rect 15215 17380 15219 17436
rect 15219 17380 15275 17436
rect 15275 17380 15279 17436
rect 15215 17376 15279 17380
rect 2861 16892 2925 16896
rect 2861 16836 2865 16892
rect 2865 16836 2921 16892
rect 2921 16836 2925 16892
rect 2861 16832 2925 16836
rect 2941 16892 3005 16896
rect 2941 16836 2945 16892
rect 2945 16836 3001 16892
rect 3001 16836 3005 16892
rect 2941 16832 3005 16836
rect 3021 16892 3085 16896
rect 3021 16836 3025 16892
rect 3025 16836 3081 16892
rect 3081 16836 3085 16892
rect 3021 16832 3085 16836
rect 3101 16892 3165 16896
rect 3101 16836 3105 16892
rect 3105 16836 3161 16892
rect 3161 16836 3165 16892
rect 3101 16832 3165 16836
rect 6679 16892 6743 16896
rect 6679 16836 6683 16892
rect 6683 16836 6739 16892
rect 6739 16836 6743 16892
rect 6679 16832 6743 16836
rect 6759 16892 6823 16896
rect 6759 16836 6763 16892
rect 6763 16836 6819 16892
rect 6819 16836 6823 16892
rect 6759 16832 6823 16836
rect 6839 16892 6903 16896
rect 6839 16836 6843 16892
rect 6843 16836 6899 16892
rect 6899 16836 6903 16892
rect 6839 16832 6903 16836
rect 6919 16892 6983 16896
rect 6919 16836 6923 16892
rect 6923 16836 6979 16892
rect 6979 16836 6983 16892
rect 6919 16832 6983 16836
rect 10497 16892 10561 16896
rect 10497 16836 10501 16892
rect 10501 16836 10557 16892
rect 10557 16836 10561 16892
rect 10497 16832 10561 16836
rect 10577 16892 10641 16896
rect 10577 16836 10581 16892
rect 10581 16836 10637 16892
rect 10637 16836 10641 16892
rect 10577 16832 10641 16836
rect 10657 16892 10721 16896
rect 10657 16836 10661 16892
rect 10661 16836 10717 16892
rect 10717 16836 10721 16892
rect 10657 16832 10721 16836
rect 10737 16892 10801 16896
rect 10737 16836 10741 16892
rect 10741 16836 10797 16892
rect 10797 16836 10801 16892
rect 10737 16832 10801 16836
rect 14315 16892 14379 16896
rect 14315 16836 14319 16892
rect 14319 16836 14375 16892
rect 14375 16836 14379 16892
rect 14315 16832 14379 16836
rect 14395 16892 14459 16896
rect 14395 16836 14399 16892
rect 14399 16836 14455 16892
rect 14455 16836 14459 16892
rect 14395 16832 14459 16836
rect 14475 16892 14539 16896
rect 14475 16836 14479 16892
rect 14479 16836 14535 16892
rect 14535 16836 14539 16892
rect 14475 16832 14539 16836
rect 14555 16892 14619 16896
rect 14555 16836 14559 16892
rect 14559 16836 14615 16892
rect 14615 16836 14619 16892
rect 14555 16832 14619 16836
rect 3521 16348 3585 16352
rect 3521 16292 3525 16348
rect 3525 16292 3581 16348
rect 3581 16292 3585 16348
rect 3521 16288 3585 16292
rect 3601 16348 3665 16352
rect 3601 16292 3605 16348
rect 3605 16292 3661 16348
rect 3661 16292 3665 16348
rect 3601 16288 3665 16292
rect 3681 16348 3745 16352
rect 3681 16292 3685 16348
rect 3685 16292 3741 16348
rect 3741 16292 3745 16348
rect 3681 16288 3745 16292
rect 3761 16348 3825 16352
rect 3761 16292 3765 16348
rect 3765 16292 3821 16348
rect 3821 16292 3825 16348
rect 3761 16288 3825 16292
rect 7339 16348 7403 16352
rect 7339 16292 7343 16348
rect 7343 16292 7399 16348
rect 7399 16292 7403 16348
rect 7339 16288 7403 16292
rect 7419 16348 7483 16352
rect 7419 16292 7423 16348
rect 7423 16292 7479 16348
rect 7479 16292 7483 16348
rect 7419 16288 7483 16292
rect 7499 16348 7563 16352
rect 7499 16292 7503 16348
rect 7503 16292 7559 16348
rect 7559 16292 7563 16348
rect 7499 16288 7563 16292
rect 7579 16348 7643 16352
rect 7579 16292 7583 16348
rect 7583 16292 7639 16348
rect 7639 16292 7643 16348
rect 7579 16288 7643 16292
rect 11157 16348 11221 16352
rect 11157 16292 11161 16348
rect 11161 16292 11217 16348
rect 11217 16292 11221 16348
rect 11157 16288 11221 16292
rect 11237 16348 11301 16352
rect 11237 16292 11241 16348
rect 11241 16292 11297 16348
rect 11297 16292 11301 16348
rect 11237 16288 11301 16292
rect 11317 16348 11381 16352
rect 11317 16292 11321 16348
rect 11321 16292 11377 16348
rect 11377 16292 11381 16348
rect 11317 16288 11381 16292
rect 11397 16348 11461 16352
rect 11397 16292 11401 16348
rect 11401 16292 11457 16348
rect 11457 16292 11461 16348
rect 11397 16288 11461 16292
rect 14975 16348 15039 16352
rect 14975 16292 14979 16348
rect 14979 16292 15035 16348
rect 15035 16292 15039 16348
rect 14975 16288 15039 16292
rect 15055 16348 15119 16352
rect 15055 16292 15059 16348
rect 15059 16292 15115 16348
rect 15115 16292 15119 16348
rect 15055 16288 15119 16292
rect 15135 16348 15199 16352
rect 15135 16292 15139 16348
rect 15139 16292 15195 16348
rect 15195 16292 15199 16348
rect 15135 16288 15199 16292
rect 15215 16348 15279 16352
rect 15215 16292 15219 16348
rect 15219 16292 15275 16348
rect 15275 16292 15279 16348
rect 15215 16288 15279 16292
rect 2861 15804 2925 15808
rect 2861 15748 2865 15804
rect 2865 15748 2921 15804
rect 2921 15748 2925 15804
rect 2861 15744 2925 15748
rect 2941 15804 3005 15808
rect 2941 15748 2945 15804
rect 2945 15748 3001 15804
rect 3001 15748 3005 15804
rect 2941 15744 3005 15748
rect 3021 15804 3085 15808
rect 3021 15748 3025 15804
rect 3025 15748 3081 15804
rect 3081 15748 3085 15804
rect 3021 15744 3085 15748
rect 3101 15804 3165 15808
rect 3101 15748 3105 15804
rect 3105 15748 3161 15804
rect 3161 15748 3165 15804
rect 3101 15744 3165 15748
rect 6679 15804 6743 15808
rect 6679 15748 6683 15804
rect 6683 15748 6739 15804
rect 6739 15748 6743 15804
rect 6679 15744 6743 15748
rect 6759 15804 6823 15808
rect 6759 15748 6763 15804
rect 6763 15748 6819 15804
rect 6819 15748 6823 15804
rect 6759 15744 6823 15748
rect 6839 15804 6903 15808
rect 6839 15748 6843 15804
rect 6843 15748 6899 15804
rect 6899 15748 6903 15804
rect 6839 15744 6903 15748
rect 6919 15804 6983 15808
rect 6919 15748 6923 15804
rect 6923 15748 6979 15804
rect 6979 15748 6983 15804
rect 6919 15744 6983 15748
rect 10497 15804 10561 15808
rect 10497 15748 10501 15804
rect 10501 15748 10557 15804
rect 10557 15748 10561 15804
rect 10497 15744 10561 15748
rect 10577 15804 10641 15808
rect 10577 15748 10581 15804
rect 10581 15748 10637 15804
rect 10637 15748 10641 15804
rect 10577 15744 10641 15748
rect 10657 15804 10721 15808
rect 10657 15748 10661 15804
rect 10661 15748 10717 15804
rect 10717 15748 10721 15804
rect 10657 15744 10721 15748
rect 10737 15804 10801 15808
rect 10737 15748 10741 15804
rect 10741 15748 10797 15804
rect 10797 15748 10801 15804
rect 10737 15744 10801 15748
rect 14315 15804 14379 15808
rect 14315 15748 14319 15804
rect 14319 15748 14375 15804
rect 14375 15748 14379 15804
rect 14315 15744 14379 15748
rect 14395 15804 14459 15808
rect 14395 15748 14399 15804
rect 14399 15748 14455 15804
rect 14455 15748 14459 15804
rect 14395 15744 14459 15748
rect 14475 15804 14539 15808
rect 14475 15748 14479 15804
rect 14479 15748 14535 15804
rect 14535 15748 14539 15804
rect 14475 15744 14539 15748
rect 14555 15804 14619 15808
rect 14555 15748 14559 15804
rect 14559 15748 14615 15804
rect 14615 15748 14619 15804
rect 14555 15744 14619 15748
rect 3521 15260 3585 15264
rect 3521 15204 3525 15260
rect 3525 15204 3581 15260
rect 3581 15204 3585 15260
rect 3521 15200 3585 15204
rect 3601 15260 3665 15264
rect 3601 15204 3605 15260
rect 3605 15204 3661 15260
rect 3661 15204 3665 15260
rect 3601 15200 3665 15204
rect 3681 15260 3745 15264
rect 3681 15204 3685 15260
rect 3685 15204 3741 15260
rect 3741 15204 3745 15260
rect 3681 15200 3745 15204
rect 3761 15260 3825 15264
rect 3761 15204 3765 15260
rect 3765 15204 3821 15260
rect 3821 15204 3825 15260
rect 3761 15200 3825 15204
rect 7339 15260 7403 15264
rect 7339 15204 7343 15260
rect 7343 15204 7399 15260
rect 7399 15204 7403 15260
rect 7339 15200 7403 15204
rect 7419 15260 7483 15264
rect 7419 15204 7423 15260
rect 7423 15204 7479 15260
rect 7479 15204 7483 15260
rect 7419 15200 7483 15204
rect 7499 15260 7563 15264
rect 7499 15204 7503 15260
rect 7503 15204 7559 15260
rect 7559 15204 7563 15260
rect 7499 15200 7563 15204
rect 7579 15260 7643 15264
rect 7579 15204 7583 15260
rect 7583 15204 7639 15260
rect 7639 15204 7643 15260
rect 7579 15200 7643 15204
rect 11157 15260 11221 15264
rect 11157 15204 11161 15260
rect 11161 15204 11217 15260
rect 11217 15204 11221 15260
rect 11157 15200 11221 15204
rect 11237 15260 11301 15264
rect 11237 15204 11241 15260
rect 11241 15204 11297 15260
rect 11297 15204 11301 15260
rect 11237 15200 11301 15204
rect 11317 15260 11381 15264
rect 11317 15204 11321 15260
rect 11321 15204 11377 15260
rect 11377 15204 11381 15260
rect 11317 15200 11381 15204
rect 11397 15260 11461 15264
rect 11397 15204 11401 15260
rect 11401 15204 11457 15260
rect 11457 15204 11461 15260
rect 11397 15200 11461 15204
rect 14975 15260 15039 15264
rect 14975 15204 14979 15260
rect 14979 15204 15035 15260
rect 15035 15204 15039 15260
rect 14975 15200 15039 15204
rect 15055 15260 15119 15264
rect 15055 15204 15059 15260
rect 15059 15204 15115 15260
rect 15115 15204 15119 15260
rect 15055 15200 15119 15204
rect 15135 15260 15199 15264
rect 15135 15204 15139 15260
rect 15139 15204 15195 15260
rect 15195 15204 15199 15260
rect 15135 15200 15199 15204
rect 15215 15260 15279 15264
rect 15215 15204 15219 15260
rect 15219 15204 15275 15260
rect 15275 15204 15279 15260
rect 15215 15200 15279 15204
rect 2861 14716 2925 14720
rect 2861 14660 2865 14716
rect 2865 14660 2921 14716
rect 2921 14660 2925 14716
rect 2861 14656 2925 14660
rect 2941 14716 3005 14720
rect 2941 14660 2945 14716
rect 2945 14660 3001 14716
rect 3001 14660 3005 14716
rect 2941 14656 3005 14660
rect 3021 14716 3085 14720
rect 3021 14660 3025 14716
rect 3025 14660 3081 14716
rect 3081 14660 3085 14716
rect 3021 14656 3085 14660
rect 3101 14716 3165 14720
rect 3101 14660 3105 14716
rect 3105 14660 3161 14716
rect 3161 14660 3165 14716
rect 3101 14656 3165 14660
rect 6679 14716 6743 14720
rect 6679 14660 6683 14716
rect 6683 14660 6739 14716
rect 6739 14660 6743 14716
rect 6679 14656 6743 14660
rect 6759 14716 6823 14720
rect 6759 14660 6763 14716
rect 6763 14660 6819 14716
rect 6819 14660 6823 14716
rect 6759 14656 6823 14660
rect 6839 14716 6903 14720
rect 6839 14660 6843 14716
rect 6843 14660 6899 14716
rect 6899 14660 6903 14716
rect 6839 14656 6903 14660
rect 6919 14716 6983 14720
rect 6919 14660 6923 14716
rect 6923 14660 6979 14716
rect 6979 14660 6983 14716
rect 6919 14656 6983 14660
rect 10497 14716 10561 14720
rect 10497 14660 10501 14716
rect 10501 14660 10557 14716
rect 10557 14660 10561 14716
rect 10497 14656 10561 14660
rect 10577 14716 10641 14720
rect 10577 14660 10581 14716
rect 10581 14660 10637 14716
rect 10637 14660 10641 14716
rect 10577 14656 10641 14660
rect 10657 14716 10721 14720
rect 10657 14660 10661 14716
rect 10661 14660 10717 14716
rect 10717 14660 10721 14716
rect 10657 14656 10721 14660
rect 10737 14716 10801 14720
rect 10737 14660 10741 14716
rect 10741 14660 10797 14716
rect 10797 14660 10801 14716
rect 10737 14656 10801 14660
rect 14315 14716 14379 14720
rect 14315 14660 14319 14716
rect 14319 14660 14375 14716
rect 14375 14660 14379 14716
rect 14315 14656 14379 14660
rect 14395 14716 14459 14720
rect 14395 14660 14399 14716
rect 14399 14660 14455 14716
rect 14455 14660 14459 14716
rect 14395 14656 14459 14660
rect 14475 14716 14539 14720
rect 14475 14660 14479 14716
rect 14479 14660 14535 14716
rect 14535 14660 14539 14716
rect 14475 14656 14539 14660
rect 14555 14716 14619 14720
rect 14555 14660 14559 14716
rect 14559 14660 14615 14716
rect 14615 14660 14619 14716
rect 14555 14656 14619 14660
rect 3521 14172 3585 14176
rect 3521 14116 3525 14172
rect 3525 14116 3581 14172
rect 3581 14116 3585 14172
rect 3521 14112 3585 14116
rect 3601 14172 3665 14176
rect 3601 14116 3605 14172
rect 3605 14116 3661 14172
rect 3661 14116 3665 14172
rect 3601 14112 3665 14116
rect 3681 14172 3745 14176
rect 3681 14116 3685 14172
rect 3685 14116 3741 14172
rect 3741 14116 3745 14172
rect 3681 14112 3745 14116
rect 3761 14172 3825 14176
rect 3761 14116 3765 14172
rect 3765 14116 3821 14172
rect 3821 14116 3825 14172
rect 3761 14112 3825 14116
rect 7339 14172 7403 14176
rect 7339 14116 7343 14172
rect 7343 14116 7399 14172
rect 7399 14116 7403 14172
rect 7339 14112 7403 14116
rect 7419 14172 7483 14176
rect 7419 14116 7423 14172
rect 7423 14116 7479 14172
rect 7479 14116 7483 14172
rect 7419 14112 7483 14116
rect 7499 14172 7563 14176
rect 7499 14116 7503 14172
rect 7503 14116 7559 14172
rect 7559 14116 7563 14172
rect 7499 14112 7563 14116
rect 7579 14172 7643 14176
rect 7579 14116 7583 14172
rect 7583 14116 7639 14172
rect 7639 14116 7643 14172
rect 7579 14112 7643 14116
rect 11157 14172 11221 14176
rect 11157 14116 11161 14172
rect 11161 14116 11217 14172
rect 11217 14116 11221 14172
rect 11157 14112 11221 14116
rect 11237 14172 11301 14176
rect 11237 14116 11241 14172
rect 11241 14116 11297 14172
rect 11297 14116 11301 14172
rect 11237 14112 11301 14116
rect 11317 14172 11381 14176
rect 11317 14116 11321 14172
rect 11321 14116 11377 14172
rect 11377 14116 11381 14172
rect 11317 14112 11381 14116
rect 11397 14172 11461 14176
rect 11397 14116 11401 14172
rect 11401 14116 11457 14172
rect 11457 14116 11461 14172
rect 11397 14112 11461 14116
rect 14975 14172 15039 14176
rect 14975 14116 14979 14172
rect 14979 14116 15035 14172
rect 15035 14116 15039 14172
rect 14975 14112 15039 14116
rect 15055 14172 15119 14176
rect 15055 14116 15059 14172
rect 15059 14116 15115 14172
rect 15115 14116 15119 14172
rect 15055 14112 15119 14116
rect 15135 14172 15199 14176
rect 15135 14116 15139 14172
rect 15139 14116 15195 14172
rect 15195 14116 15199 14172
rect 15135 14112 15199 14116
rect 15215 14172 15279 14176
rect 15215 14116 15219 14172
rect 15219 14116 15275 14172
rect 15275 14116 15279 14172
rect 15215 14112 15279 14116
rect 2861 13628 2925 13632
rect 2861 13572 2865 13628
rect 2865 13572 2921 13628
rect 2921 13572 2925 13628
rect 2861 13568 2925 13572
rect 2941 13628 3005 13632
rect 2941 13572 2945 13628
rect 2945 13572 3001 13628
rect 3001 13572 3005 13628
rect 2941 13568 3005 13572
rect 3021 13628 3085 13632
rect 3021 13572 3025 13628
rect 3025 13572 3081 13628
rect 3081 13572 3085 13628
rect 3021 13568 3085 13572
rect 3101 13628 3165 13632
rect 3101 13572 3105 13628
rect 3105 13572 3161 13628
rect 3161 13572 3165 13628
rect 3101 13568 3165 13572
rect 6679 13628 6743 13632
rect 6679 13572 6683 13628
rect 6683 13572 6739 13628
rect 6739 13572 6743 13628
rect 6679 13568 6743 13572
rect 6759 13628 6823 13632
rect 6759 13572 6763 13628
rect 6763 13572 6819 13628
rect 6819 13572 6823 13628
rect 6759 13568 6823 13572
rect 6839 13628 6903 13632
rect 6839 13572 6843 13628
rect 6843 13572 6899 13628
rect 6899 13572 6903 13628
rect 6839 13568 6903 13572
rect 6919 13628 6983 13632
rect 6919 13572 6923 13628
rect 6923 13572 6979 13628
rect 6979 13572 6983 13628
rect 6919 13568 6983 13572
rect 10497 13628 10561 13632
rect 10497 13572 10501 13628
rect 10501 13572 10557 13628
rect 10557 13572 10561 13628
rect 10497 13568 10561 13572
rect 10577 13628 10641 13632
rect 10577 13572 10581 13628
rect 10581 13572 10637 13628
rect 10637 13572 10641 13628
rect 10577 13568 10641 13572
rect 10657 13628 10721 13632
rect 10657 13572 10661 13628
rect 10661 13572 10717 13628
rect 10717 13572 10721 13628
rect 10657 13568 10721 13572
rect 10737 13628 10801 13632
rect 10737 13572 10741 13628
rect 10741 13572 10797 13628
rect 10797 13572 10801 13628
rect 10737 13568 10801 13572
rect 14315 13628 14379 13632
rect 14315 13572 14319 13628
rect 14319 13572 14375 13628
rect 14375 13572 14379 13628
rect 14315 13568 14379 13572
rect 14395 13628 14459 13632
rect 14395 13572 14399 13628
rect 14399 13572 14455 13628
rect 14455 13572 14459 13628
rect 14395 13568 14459 13572
rect 14475 13628 14539 13632
rect 14475 13572 14479 13628
rect 14479 13572 14535 13628
rect 14535 13572 14539 13628
rect 14475 13568 14539 13572
rect 14555 13628 14619 13632
rect 14555 13572 14559 13628
rect 14559 13572 14615 13628
rect 14615 13572 14619 13628
rect 14555 13568 14619 13572
rect 3521 13084 3585 13088
rect 3521 13028 3525 13084
rect 3525 13028 3581 13084
rect 3581 13028 3585 13084
rect 3521 13024 3585 13028
rect 3601 13084 3665 13088
rect 3601 13028 3605 13084
rect 3605 13028 3661 13084
rect 3661 13028 3665 13084
rect 3601 13024 3665 13028
rect 3681 13084 3745 13088
rect 3681 13028 3685 13084
rect 3685 13028 3741 13084
rect 3741 13028 3745 13084
rect 3681 13024 3745 13028
rect 3761 13084 3825 13088
rect 3761 13028 3765 13084
rect 3765 13028 3821 13084
rect 3821 13028 3825 13084
rect 3761 13024 3825 13028
rect 7339 13084 7403 13088
rect 7339 13028 7343 13084
rect 7343 13028 7399 13084
rect 7399 13028 7403 13084
rect 7339 13024 7403 13028
rect 7419 13084 7483 13088
rect 7419 13028 7423 13084
rect 7423 13028 7479 13084
rect 7479 13028 7483 13084
rect 7419 13024 7483 13028
rect 7499 13084 7563 13088
rect 7499 13028 7503 13084
rect 7503 13028 7559 13084
rect 7559 13028 7563 13084
rect 7499 13024 7563 13028
rect 7579 13084 7643 13088
rect 7579 13028 7583 13084
rect 7583 13028 7639 13084
rect 7639 13028 7643 13084
rect 7579 13024 7643 13028
rect 11157 13084 11221 13088
rect 11157 13028 11161 13084
rect 11161 13028 11217 13084
rect 11217 13028 11221 13084
rect 11157 13024 11221 13028
rect 11237 13084 11301 13088
rect 11237 13028 11241 13084
rect 11241 13028 11297 13084
rect 11297 13028 11301 13084
rect 11237 13024 11301 13028
rect 11317 13084 11381 13088
rect 11317 13028 11321 13084
rect 11321 13028 11377 13084
rect 11377 13028 11381 13084
rect 11317 13024 11381 13028
rect 11397 13084 11461 13088
rect 11397 13028 11401 13084
rect 11401 13028 11457 13084
rect 11457 13028 11461 13084
rect 11397 13024 11461 13028
rect 14975 13084 15039 13088
rect 14975 13028 14979 13084
rect 14979 13028 15035 13084
rect 15035 13028 15039 13084
rect 14975 13024 15039 13028
rect 15055 13084 15119 13088
rect 15055 13028 15059 13084
rect 15059 13028 15115 13084
rect 15115 13028 15119 13084
rect 15055 13024 15119 13028
rect 15135 13084 15199 13088
rect 15135 13028 15139 13084
rect 15139 13028 15195 13084
rect 15195 13028 15199 13084
rect 15135 13024 15199 13028
rect 15215 13084 15279 13088
rect 15215 13028 15219 13084
rect 15219 13028 15275 13084
rect 15275 13028 15279 13084
rect 15215 13024 15279 13028
rect 2861 12540 2925 12544
rect 2861 12484 2865 12540
rect 2865 12484 2921 12540
rect 2921 12484 2925 12540
rect 2861 12480 2925 12484
rect 2941 12540 3005 12544
rect 2941 12484 2945 12540
rect 2945 12484 3001 12540
rect 3001 12484 3005 12540
rect 2941 12480 3005 12484
rect 3021 12540 3085 12544
rect 3021 12484 3025 12540
rect 3025 12484 3081 12540
rect 3081 12484 3085 12540
rect 3021 12480 3085 12484
rect 3101 12540 3165 12544
rect 3101 12484 3105 12540
rect 3105 12484 3161 12540
rect 3161 12484 3165 12540
rect 3101 12480 3165 12484
rect 6679 12540 6743 12544
rect 6679 12484 6683 12540
rect 6683 12484 6739 12540
rect 6739 12484 6743 12540
rect 6679 12480 6743 12484
rect 6759 12540 6823 12544
rect 6759 12484 6763 12540
rect 6763 12484 6819 12540
rect 6819 12484 6823 12540
rect 6759 12480 6823 12484
rect 6839 12540 6903 12544
rect 6839 12484 6843 12540
rect 6843 12484 6899 12540
rect 6899 12484 6903 12540
rect 6839 12480 6903 12484
rect 6919 12540 6983 12544
rect 6919 12484 6923 12540
rect 6923 12484 6979 12540
rect 6979 12484 6983 12540
rect 6919 12480 6983 12484
rect 10497 12540 10561 12544
rect 10497 12484 10501 12540
rect 10501 12484 10557 12540
rect 10557 12484 10561 12540
rect 10497 12480 10561 12484
rect 10577 12540 10641 12544
rect 10577 12484 10581 12540
rect 10581 12484 10637 12540
rect 10637 12484 10641 12540
rect 10577 12480 10641 12484
rect 10657 12540 10721 12544
rect 10657 12484 10661 12540
rect 10661 12484 10717 12540
rect 10717 12484 10721 12540
rect 10657 12480 10721 12484
rect 10737 12540 10801 12544
rect 10737 12484 10741 12540
rect 10741 12484 10797 12540
rect 10797 12484 10801 12540
rect 10737 12480 10801 12484
rect 14315 12540 14379 12544
rect 14315 12484 14319 12540
rect 14319 12484 14375 12540
rect 14375 12484 14379 12540
rect 14315 12480 14379 12484
rect 14395 12540 14459 12544
rect 14395 12484 14399 12540
rect 14399 12484 14455 12540
rect 14455 12484 14459 12540
rect 14395 12480 14459 12484
rect 14475 12540 14539 12544
rect 14475 12484 14479 12540
rect 14479 12484 14535 12540
rect 14535 12484 14539 12540
rect 14475 12480 14539 12484
rect 14555 12540 14619 12544
rect 14555 12484 14559 12540
rect 14559 12484 14615 12540
rect 14615 12484 14619 12540
rect 14555 12480 14619 12484
rect 3521 11996 3585 12000
rect 3521 11940 3525 11996
rect 3525 11940 3581 11996
rect 3581 11940 3585 11996
rect 3521 11936 3585 11940
rect 3601 11996 3665 12000
rect 3601 11940 3605 11996
rect 3605 11940 3661 11996
rect 3661 11940 3665 11996
rect 3601 11936 3665 11940
rect 3681 11996 3745 12000
rect 3681 11940 3685 11996
rect 3685 11940 3741 11996
rect 3741 11940 3745 11996
rect 3681 11936 3745 11940
rect 3761 11996 3825 12000
rect 3761 11940 3765 11996
rect 3765 11940 3821 11996
rect 3821 11940 3825 11996
rect 3761 11936 3825 11940
rect 7339 11996 7403 12000
rect 7339 11940 7343 11996
rect 7343 11940 7399 11996
rect 7399 11940 7403 11996
rect 7339 11936 7403 11940
rect 7419 11996 7483 12000
rect 7419 11940 7423 11996
rect 7423 11940 7479 11996
rect 7479 11940 7483 11996
rect 7419 11936 7483 11940
rect 7499 11996 7563 12000
rect 7499 11940 7503 11996
rect 7503 11940 7559 11996
rect 7559 11940 7563 11996
rect 7499 11936 7563 11940
rect 7579 11996 7643 12000
rect 7579 11940 7583 11996
rect 7583 11940 7639 11996
rect 7639 11940 7643 11996
rect 7579 11936 7643 11940
rect 11157 11996 11221 12000
rect 11157 11940 11161 11996
rect 11161 11940 11217 11996
rect 11217 11940 11221 11996
rect 11157 11936 11221 11940
rect 11237 11996 11301 12000
rect 11237 11940 11241 11996
rect 11241 11940 11297 11996
rect 11297 11940 11301 11996
rect 11237 11936 11301 11940
rect 11317 11996 11381 12000
rect 11317 11940 11321 11996
rect 11321 11940 11377 11996
rect 11377 11940 11381 11996
rect 11317 11936 11381 11940
rect 11397 11996 11461 12000
rect 11397 11940 11401 11996
rect 11401 11940 11457 11996
rect 11457 11940 11461 11996
rect 11397 11936 11461 11940
rect 14975 11996 15039 12000
rect 14975 11940 14979 11996
rect 14979 11940 15035 11996
rect 15035 11940 15039 11996
rect 14975 11936 15039 11940
rect 15055 11996 15119 12000
rect 15055 11940 15059 11996
rect 15059 11940 15115 11996
rect 15115 11940 15119 11996
rect 15055 11936 15119 11940
rect 15135 11996 15199 12000
rect 15135 11940 15139 11996
rect 15139 11940 15195 11996
rect 15195 11940 15199 11996
rect 15135 11936 15199 11940
rect 15215 11996 15279 12000
rect 15215 11940 15219 11996
rect 15219 11940 15275 11996
rect 15275 11940 15279 11996
rect 15215 11936 15279 11940
rect 2861 11452 2925 11456
rect 2861 11396 2865 11452
rect 2865 11396 2921 11452
rect 2921 11396 2925 11452
rect 2861 11392 2925 11396
rect 2941 11452 3005 11456
rect 2941 11396 2945 11452
rect 2945 11396 3001 11452
rect 3001 11396 3005 11452
rect 2941 11392 3005 11396
rect 3021 11452 3085 11456
rect 3021 11396 3025 11452
rect 3025 11396 3081 11452
rect 3081 11396 3085 11452
rect 3021 11392 3085 11396
rect 3101 11452 3165 11456
rect 3101 11396 3105 11452
rect 3105 11396 3161 11452
rect 3161 11396 3165 11452
rect 3101 11392 3165 11396
rect 6679 11452 6743 11456
rect 6679 11396 6683 11452
rect 6683 11396 6739 11452
rect 6739 11396 6743 11452
rect 6679 11392 6743 11396
rect 6759 11452 6823 11456
rect 6759 11396 6763 11452
rect 6763 11396 6819 11452
rect 6819 11396 6823 11452
rect 6759 11392 6823 11396
rect 6839 11452 6903 11456
rect 6839 11396 6843 11452
rect 6843 11396 6899 11452
rect 6899 11396 6903 11452
rect 6839 11392 6903 11396
rect 6919 11452 6983 11456
rect 6919 11396 6923 11452
rect 6923 11396 6979 11452
rect 6979 11396 6983 11452
rect 6919 11392 6983 11396
rect 10497 11452 10561 11456
rect 10497 11396 10501 11452
rect 10501 11396 10557 11452
rect 10557 11396 10561 11452
rect 10497 11392 10561 11396
rect 10577 11452 10641 11456
rect 10577 11396 10581 11452
rect 10581 11396 10637 11452
rect 10637 11396 10641 11452
rect 10577 11392 10641 11396
rect 10657 11452 10721 11456
rect 10657 11396 10661 11452
rect 10661 11396 10717 11452
rect 10717 11396 10721 11452
rect 10657 11392 10721 11396
rect 10737 11452 10801 11456
rect 10737 11396 10741 11452
rect 10741 11396 10797 11452
rect 10797 11396 10801 11452
rect 10737 11392 10801 11396
rect 14315 11452 14379 11456
rect 14315 11396 14319 11452
rect 14319 11396 14375 11452
rect 14375 11396 14379 11452
rect 14315 11392 14379 11396
rect 14395 11452 14459 11456
rect 14395 11396 14399 11452
rect 14399 11396 14455 11452
rect 14455 11396 14459 11452
rect 14395 11392 14459 11396
rect 14475 11452 14539 11456
rect 14475 11396 14479 11452
rect 14479 11396 14535 11452
rect 14535 11396 14539 11452
rect 14475 11392 14539 11396
rect 14555 11452 14619 11456
rect 14555 11396 14559 11452
rect 14559 11396 14615 11452
rect 14615 11396 14619 11452
rect 14555 11392 14619 11396
rect 3521 10908 3585 10912
rect 3521 10852 3525 10908
rect 3525 10852 3581 10908
rect 3581 10852 3585 10908
rect 3521 10848 3585 10852
rect 3601 10908 3665 10912
rect 3601 10852 3605 10908
rect 3605 10852 3661 10908
rect 3661 10852 3665 10908
rect 3601 10848 3665 10852
rect 3681 10908 3745 10912
rect 3681 10852 3685 10908
rect 3685 10852 3741 10908
rect 3741 10852 3745 10908
rect 3681 10848 3745 10852
rect 3761 10908 3825 10912
rect 3761 10852 3765 10908
rect 3765 10852 3821 10908
rect 3821 10852 3825 10908
rect 3761 10848 3825 10852
rect 7339 10908 7403 10912
rect 7339 10852 7343 10908
rect 7343 10852 7399 10908
rect 7399 10852 7403 10908
rect 7339 10848 7403 10852
rect 7419 10908 7483 10912
rect 7419 10852 7423 10908
rect 7423 10852 7479 10908
rect 7479 10852 7483 10908
rect 7419 10848 7483 10852
rect 7499 10908 7563 10912
rect 7499 10852 7503 10908
rect 7503 10852 7559 10908
rect 7559 10852 7563 10908
rect 7499 10848 7563 10852
rect 7579 10908 7643 10912
rect 7579 10852 7583 10908
rect 7583 10852 7639 10908
rect 7639 10852 7643 10908
rect 7579 10848 7643 10852
rect 11157 10908 11221 10912
rect 11157 10852 11161 10908
rect 11161 10852 11217 10908
rect 11217 10852 11221 10908
rect 11157 10848 11221 10852
rect 11237 10908 11301 10912
rect 11237 10852 11241 10908
rect 11241 10852 11297 10908
rect 11297 10852 11301 10908
rect 11237 10848 11301 10852
rect 11317 10908 11381 10912
rect 11317 10852 11321 10908
rect 11321 10852 11377 10908
rect 11377 10852 11381 10908
rect 11317 10848 11381 10852
rect 11397 10908 11461 10912
rect 11397 10852 11401 10908
rect 11401 10852 11457 10908
rect 11457 10852 11461 10908
rect 11397 10848 11461 10852
rect 14975 10908 15039 10912
rect 14975 10852 14979 10908
rect 14979 10852 15035 10908
rect 15035 10852 15039 10908
rect 14975 10848 15039 10852
rect 15055 10908 15119 10912
rect 15055 10852 15059 10908
rect 15059 10852 15115 10908
rect 15115 10852 15119 10908
rect 15055 10848 15119 10852
rect 15135 10908 15199 10912
rect 15135 10852 15139 10908
rect 15139 10852 15195 10908
rect 15195 10852 15199 10908
rect 15135 10848 15199 10852
rect 15215 10908 15279 10912
rect 15215 10852 15219 10908
rect 15219 10852 15275 10908
rect 15275 10852 15279 10908
rect 15215 10848 15279 10852
rect 2861 10364 2925 10368
rect 2861 10308 2865 10364
rect 2865 10308 2921 10364
rect 2921 10308 2925 10364
rect 2861 10304 2925 10308
rect 2941 10364 3005 10368
rect 2941 10308 2945 10364
rect 2945 10308 3001 10364
rect 3001 10308 3005 10364
rect 2941 10304 3005 10308
rect 3021 10364 3085 10368
rect 3021 10308 3025 10364
rect 3025 10308 3081 10364
rect 3081 10308 3085 10364
rect 3021 10304 3085 10308
rect 3101 10364 3165 10368
rect 3101 10308 3105 10364
rect 3105 10308 3161 10364
rect 3161 10308 3165 10364
rect 3101 10304 3165 10308
rect 6679 10364 6743 10368
rect 6679 10308 6683 10364
rect 6683 10308 6739 10364
rect 6739 10308 6743 10364
rect 6679 10304 6743 10308
rect 6759 10364 6823 10368
rect 6759 10308 6763 10364
rect 6763 10308 6819 10364
rect 6819 10308 6823 10364
rect 6759 10304 6823 10308
rect 6839 10364 6903 10368
rect 6839 10308 6843 10364
rect 6843 10308 6899 10364
rect 6899 10308 6903 10364
rect 6839 10304 6903 10308
rect 6919 10364 6983 10368
rect 6919 10308 6923 10364
rect 6923 10308 6979 10364
rect 6979 10308 6983 10364
rect 6919 10304 6983 10308
rect 10497 10364 10561 10368
rect 10497 10308 10501 10364
rect 10501 10308 10557 10364
rect 10557 10308 10561 10364
rect 10497 10304 10561 10308
rect 10577 10364 10641 10368
rect 10577 10308 10581 10364
rect 10581 10308 10637 10364
rect 10637 10308 10641 10364
rect 10577 10304 10641 10308
rect 10657 10364 10721 10368
rect 10657 10308 10661 10364
rect 10661 10308 10717 10364
rect 10717 10308 10721 10364
rect 10657 10304 10721 10308
rect 10737 10364 10801 10368
rect 10737 10308 10741 10364
rect 10741 10308 10797 10364
rect 10797 10308 10801 10364
rect 10737 10304 10801 10308
rect 14315 10364 14379 10368
rect 14315 10308 14319 10364
rect 14319 10308 14375 10364
rect 14375 10308 14379 10364
rect 14315 10304 14379 10308
rect 14395 10364 14459 10368
rect 14395 10308 14399 10364
rect 14399 10308 14455 10364
rect 14455 10308 14459 10364
rect 14395 10304 14459 10308
rect 14475 10364 14539 10368
rect 14475 10308 14479 10364
rect 14479 10308 14535 10364
rect 14535 10308 14539 10364
rect 14475 10304 14539 10308
rect 14555 10364 14619 10368
rect 14555 10308 14559 10364
rect 14559 10308 14615 10364
rect 14615 10308 14619 10364
rect 14555 10304 14619 10308
rect 3521 9820 3585 9824
rect 3521 9764 3525 9820
rect 3525 9764 3581 9820
rect 3581 9764 3585 9820
rect 3521 9760 3585 9764
rect 3601 9820 3665 9824
rect 3601 9764 3605 9820
rect 3605 9764 3661 9820
rect 3661 9764 3665 9820
rect 3601 9760 3665 9764
rect 3681 9820 3745 9824
rect 3681 9764 3685 9820
rect 3685 9764 3741 9820
rect 3741 9764 3745 9820
rect 3681 9760 3745 9764
rect 3761 9820 3825 9824
rect 3761 9764 3765 9820
rect 3765 9764 3821 9820
rect 3821 9764 3825 9820
rect 3761 9760 3825 9764
rect 7339 9820 7403 9824
rect 7339 9764 7343 9820
rect 7343 9764 7399 9820
rect 7399 9764 7403 9820
rect 7339 9760 7403 9764
rect 7419 9820 7483 9824
rect 7419 9764 7423 9820
rect 7423 9764 7479 9820
rect 7479 9764 7483 9820
rect 7419 9760 7483 9764
rect 7499 9820 7563 9824
rect 7499 9764 7503 9820
rect 7503 9764 7559 9820
rect 7559 9764 7563 9820
rect 7499 9760 7563 9764
rect 7579 9820 7643 9824
rect 7579 9764 7583 9820
rect 7583 9764 7639 9820
rect 7639 9764 7643 9820
rect 7579 9760 7643 9764
rect 11157 9820 11221 9824
rect 11157 9764 11161 9820
rect 11161 9764 11217 9820
rect 11217 9764 11221 9820
rect 11157 9760 11221 9764
rect 11237 9820 11301 9824
rect 11237 9764 11241 9820
rect 11241 9764 11297 9820
rect 11297 9764 11301 9820
rect 11237 9760 11301 9764
rect 11317 9820 11381 9824
rect 11317 9764 11321 9820
rect 11321 9764 11377 9820
rect 11377 9764 11381 9820
rect 11317 9760 11381 9764
rect 11397 9820 11461 9824
rect 11397 9764 11401 9820
rect 11401 9764 11457 9820
rect 11457 9764 11461 9820
rect 11397 9760 11461 9764
rect 14975 9820 15039 9824
rect 14975 9764 14979 9820
rect 14979 9764 15035 9820
rect 15035 9764 15039 9820
rect 14975 9760 15039 9764
rect 15055 9820 15119 9824
rect 15055 9764 15059 9820
rect 15059 9764 15115 9820
rect 15115 9764 15119 9820
rect 15055 9760 15119 9764
rect 15135 9820 15199 9824
rect 15135 9764 15139 9820
rect 15139 9764 15195 9820
rect 15195 9764 15199 9820
rect 15135 9760 15199 9764
rect 15215 9820 15279 9824
rect 15215 9764 15219 9820
rect 15219 9764 15275 9820
rect 15275 9764 15279 9820
rect 15215 9760 15279 9764
rect 2861 9276 2925 9280
rect 2861 9220 2865 9276
rect 2865 9220 2921 9276
rect 2921 9220 2925 9276
rect 2861 9216 2925 9220
rect 2941 9276 3005 9280
rect 2941 9220 2945 9276
rect 2945 9220 3001 9276
rect 3001 9220 3005 9276
rect 2941 9216 3005 9220
rect 3021 9276 3085 9280
rect 3021 9220 3025 9276
rect 3025 9220 3081 9276
rect 3081 9220 3085 9276
rect 3021 9216 3085 9220
rect 3101 9276 3165 9280
rect 3101 9220 3105 9276
rect 3105 9220 3161 9276
rect 3161 9220 3165 9276
rect 3101 9216 3165 9220
rect 6679 9276 6743 9280
rect 6679 9220 6683 9276
rect 6683 9220 6739 9276
rect 6739 9220 6743 9276
rect 6679 9216 6743 9220
rect 6759 9276 6823 9280
rect 6759 9220 6763 9276
rect 6763 9220 6819 9276
rect 6819 9220 6823 9276
rect 6759 9216 6823 9220
rect 6839 9276 6903 9280
rect 6839 9220 6843 9276
rect 6843 9220 6899 9276
rect 6899 9220 6903 9276
rect 6839 9216 6903 9220
rect 6919 9276 6983 9280
rect 6919 9220 6923 9276
rect 6923 9220 6979 9276
rect 6979 9220 6983 9276
rect 6919 9216 6983 9220
rect 10497 9276 10561 9280
rect 10497 9220 10501 9276
rect 10501 9220 10557 9276
rect 10557 9220 10561 9276
rect 10497 9216 10561 9220
rect 10577 9276 10641 9280
rect 10577 9220 10581 9276
rect 10581 9220 10637 9276
rect 10637 9220 10641 9276
rect 10577 9216 10641 9220
rect 10657 9276 10721 9280
rect 10657 9220 10661 9276
rect 10661 9220 10717 9276
rect 10717 9220 10721 9276
rect 10657 9216 10721 9220
rect 10737 9276 10801 9280
rect 10737 9220 10741 9276
rect 10741 9220 10797 9276
rect 10797 9220 10801 9276
rect 10737 9216 10801 9220
rect 14315 9276 14379 9280
rect 14315 9220 14319 9276
rect 14319 9220 14375 9276
rect 14375 9220 14379 9276
rect 14315 9216 14379 9220
rect 14395 9276 14459 9280
rect 14395 9220 14399 9276
rect 14399 9220 14455 9276
rect 14455 9220 14459 9276
rect 14395 9216 14459 9220
rect 14475 9276 14539 9280
rect 14475 9220 14479 9276
rect 14479 9220 14535 9276
rect 14535 9220 14539 9276
rect 14475 9216 14539 9220
rect 14555 9276 14619 9280
rect 14555 9220 14559 9276
rect 14559 9220 14615 9276
rect 14615 9220 14619 9276
rect 14555 9216 14619 9220
rect 3521 8732 3585 8736
rect 3521 8676 3525 8732
rect 3525 8676 3581 8732
rect 3581 8676 3585 8732
rect 3521 8672 3585 8676
rect 3601 8732 3665 8736
rect 3601 8676 3605 8732
rect 3605 8676 3661 8732
rect 3661 8676 3665 8732
rect 3601 8672 3665 8676
rect 3681 8732 3745 8736
rect 3681 8676 3685 8732
rect 3685 8676 3741 8732
rect 3741 8676 3745 8732
rect 3681 8672 3745 8676
rect 3761 8732 3825 8736
rect 3761 8676 3765 8732
rect 3765 8676 3821 8732
rect 3821 8676 3825 8732
rect 3761 8672 3825 8676
rect 7339 8732 7403 8736
rect 7339 8676 7343 8732
rect 7343 8676 7399 8732
rect 7399 8676 7403 8732
rect 7339 8672 7403 8676
rect 7419 8732 7483 8736
rect 7419 8676 7423 8732
rect 7423 8676 7479 8732
rect 7479 8676 7483 8732
rect 7419 8672 7483 8676
rect 7499 8732 7563 8736
rect 7499 8676 7503 8732
rect 7503 8676 7559 8732
rect 7559 8676 7563 8732
rect 7499 8672 7563 8676
rect 7579 8732 7643 8736
rect 7579 8676 7583 8732
rect 7583 8676 7639 8732
rect 7639 8676 7643 8732
rect 7579 8672 7643 8676
rect 11157 8732 11221 8736
rect 11157 8676 11161 8732
rect 11161 8676 11217 8732
rect 11217 8676 11221 8732
rect 11157 8672 11221 8676
rect 11237 8732 11301 8736
rect 11237 8676 11241 8732
rect 11241 8676 11297 8732
rect 11297 8676 11301 8732
rect 11237 8672 11301 8676
rect 11317 8732 11381 8736
rect 11317 8676 11321 8732
rect 11321 8676 11377 8732
rect 11377 8676 11381 8732
rect 11317 8672 11381 8676
rect 11397 8732 11461 8736
rect 11397 8676 11401 8732
rect 11401 8676 11457 8732
rect 11457 8676 11461 8732
rect 11397 8672 11461 8676
rect 14975 8732 15039 8736
rect 14975 8676 14979 8732
rect 14979 8676 15035 8732
rect 15035 8676 15039 8732
rect 14975 8672 15039 8676
rect 15055 8732 15119 8736
rect 15055 8676 15059 8732
rect 15059 8676 15115 8732
rect 15115 8676 15119 8732
rect 15055 8672 15119 8676
rect 15135 8732 15199 8736
rect 15135 8676 15139 8732
rect 15139 8676 15195 8732
rect 15195 8676 15199 8732
rect 15135 8672 15199 8676
rect 15215 8732 15279 8736
rect 15215 8676 15219 8732
rect 15219 8676 15275 8732
rect 15275 8676 15279 8732
rect 15215 8672 15279 8676
rect 2861 8188 2925 8192
rect 2861 8132 2865 8188
rect 2865 8132 2921 8188
rect 2921 8132 2925 8188
rect 2861 8128 2925 8132
rect 2941 8188 3005 8192
rect 2941 8132 2945 8188
rect 2945 8132 3001 8188
rect 3001 8132 3005 8188
rect 2941 8128 3005 8132
rect 3021 8188 3085 8192
rect 3021 8132 3025 8188
rect 3025 8132 3081 8188
rect 3081 8132 3085 8188
rect 3021 8128 3085 8132
rect 3101 8188 3165 8192
rect 3101 8132 3105 8188
rect 3105 8132 3161 8188
rect 3161 8132 3165 8188
rect 3101 8128 3165 8132
rect 6679 8188 6743 8192
rect 6679 8132 6683 8188
rect 6683 8132 6739 8188
rect 6739 8132 6743 8188
rect 6679 8128 6743 8132
rect 6759 8188 6823 8192
rect 6759 8132 6763 8188
rect 6763 8132 6819 8188
rect 6819 8132 6823 8188
rect 6759 8128 6823 8132
rect 6839 8188 6903 8192
rect 6839 8132 6843 8188
rect 6843 8132 6899 8188
rect 6899 8132 6903 8188
rect 6839 8128 6903 8132
rect 6919 8188 6983 8192
rect 6919 8132 6923 8188
rect 6923 8132 6979 8188
rect 6979 8132 6983 8188
rect 6919 8128 6983 8132
rect 10497 8188 10561 8192
rect 10497 8132 10501 8188
rect 10501 8132 10557 8188
rect 10557 8132 10561 8188
rect 10497 8128 10561 8132
rect 10577 8188 10641 8192
rect 10577 8132 10581 8188
rect 10581 8132 10637 8188
rect 10637 8132 10641 8188
rect 10577 8128 10641 8132
rect 10657 8188 10721 8192
rect 10657 8132 10661 8188
rect 10661 8132 10717 8188
rect 10717 8132 10721 8188
rect 10657 8128 10721 8132
rect 10737 8188 10801 8192
rect 10737 8132 10741 8188
rect 10741 8132 10797 8188
rect 10797 8132 10801 8188
rect 10737 8128 10801 8132
rect 14315 8188 14379 8192
rect 14315 8132 14319 8188
rect 14319 8132 14375 8188
rect 14375 8132 14379 8188
rect 14315 8128 14379 8132
rect 14395 8188 14459 8192
rect 14395 8132 14399 8188
rect 14399 8132 14455 8188
rect 14455 8132 14459 8188
rect 14395 8128 14459 8132
rect 14475 8188 14539 8192
rect 14475 8132 14479 8188
rect 14479 8132 14535 8188
rect 14535 8132 14539 8188
rect 14475 8128 14539 8132
rect 14555 8188 14619 8192
rect 14555 8132 14559 8188
rect 14559 8132 14615 8188
rect 14615 8132 14619 8188
rect 14555 8128 14619 8132
rect 3521 7644 3585 7648
rect 3521 7588 3525 7644
rect 3525 7588 3581 7644
rect 3581 7588 3585 7644
rect 3521 7584 3585 7588
rect 3601 7644 3665 7648
rect 3601 7588 3605 7644
rect 3605 7588 3661 7644
rect 3661 7588 3665 7644
rect 3601 7584 3665 7588
rect 3681 7644 3745 7648
rect 3681 7588 3685 7644
rect 3685 7588 3741 7644
rect 3741 7588 3745 7644
rect 3681 7584 3745 7588
rect 3761 7644 3825 7648
rect 3761 7588 3765 7644
rect 3765 7588 3821 7644
rect 3821 7588 3825 7644
rect 3761 7584 3825 7588
rect 7339 7644 7403 7648
rect 7339 7588 7343 7644
rect 7343 7588 7399 7644
rect 7399 7588 7403 7644
rect 7339 7584 7403 7588
rect 7419 7644 7483 7648
rect 7419 7588 7423 7644
rect 7423 7588 7479 7644
rect 7479 7588 7483 7644
rect 7419 7584 7483 7588
rect 7499 7644 7563 7648
rect 7499 7588 7503 7644
rect 7503 7588 7559 7644
rect 7559 7588 7563 7644
rect 7499 7584 7563 7588
rect 7579 7644 7643 7648
rect 7579 7588 7583 7644
rect 7583 7588 7639 7644
rect 7639 7588 7643 7644
rect 7579 7584 7643 7588
rect 11157 7644 11221 7648
rect 11157 7588 11161 7644
rect 11161 7588 11217 7644
rect 11217 7588 11221 7644
rect 11157 7584 11221 7588
rect 11237 7644 11301 7648
rect 11237 7588 11241 7644
rect 11241 7588 11297 7644
rect 11297 7588 11301 7644
rect 11237 7584 11301 7588
rect 11317 7644 11381 7648
rect 11317 7588 11321 7644
rect 11321 7588 11377 7644
rect 11377 7588 11381 7644
rect 11317 7584 11381 7588
rect 11397 7644 11461 7648
rect 11397 7588 11401 7644
rect 11401 7588 11457 7644
rect 11457 7588 11461 7644
rect 11397 7584 11461 7588
rect 14975 7644 15039 7648
rect 14975 7588 14979 7644
rect 14979 7588 15035 7644
rect 15035 7588 15039 7644
rect 14975 7584 15039 7588
rect 15055 7644 15119 7648
rect 15055 7588 15059 7644
rect 15059 7588 15115 7644
rect 15115 7588 15119 7644
rect 15055 7584 15119 7588
rect 15135 7644 15199 7648
rect 15135 7588 15139 7644
rect 15139 7588 15195 7644
rect 15195 7588 15199 7644
rect 15135 7584 15199 7588
rect 15215 7644 15279 7648
rect 15215 7588 15219 7644
rect 15219 7588 15275 7644
rect 15275 7588 15279 7644
rect 15215 7584 15279 7588
rect 2861 7100 2925 7104
rect 2861 7044 2865 7100
rect 2865 7044 2921 7100
rect 2921 7044 2925 7100
rect 2861 7040 2925 7044
rect 2941 7100 3005 7104
rect 2941 7044 2945 7100
rect 2945 7044 3001 7100
rect 3001 7044 3005 7100
rect 2941 7040 3005 7044
rect 3021 7100 3085 7104
rect 3021 7044 3025 7100
rect 3025 7044 3081 7100
rect 3081 7044 3085 7100
rect 3021 7040 3085 7044
rect 3101 7100 3165 7104
rect 3101 7044 3105 7100
rect 3105 7044 3161 7100
rect 3161 7044 3165 7100
rect 3101 7040 3165 7044
rect 6679 7100 6743 7104
rect 6679 7044 6683 7100
rect 6683 7044 6739 7100
rect 6739 7044 6743 7100
rect 6679 7040 6743 7044
rect 6759 7100 6823 7104
rect 6759 7044 6763 7100
rect 6763 7044 6819 7100
rect 6819 7044 6823 7100
rect 6759 7040 6823 7044
rect 6839 7100 6903 7104
rect 6839 7044 6843 7100
rect 6843 7044 6899 7100
rect 6899 7044 6903 7100
rect 6839 7040 6903 7044
rect 6919 7100 6983 7104
rect 6919 7044 6923 7100
rect 6923 7044 6979 7100
rect 6979 7044 6983 7100
rect 6919 7040 6983 7044
rect 10497 7100 10561 7104
rect 10497 7044 10501 7100
rect 10501 7044 10557 7100
rect 10557 7044 10561 7100
rect 10497 7040 10561 7044
rect 10577 7100 10641 7104
rect 10577 7044 10581 7100
rect 10581 7044 10637 7100
rect 10637 7044 10641 7100
rect 10577 7040 10641 7044
rect 10657 7100 10721 7104
rect 10657 7044 10661 7100
rect 10661 7044 10717 7100
rect 10717 7044 10721 7100
rect 10657 7040 10721 7044
rect 10737 7100 10801 7104
rect 10737 7044 10741 7100
rect 10741 7044 10797 7100
rect 10797 7044 10801 7100
rect 10737 7040 10801 7044
rect 14315 7100 14379 7104
rect 14315 7044 14319 7100
rect 14319 7044 14375 7100
rect 14375 7044 14379 7100
rect 14315 7040 14379 7044
rect 14395 7100 14459 7104
rect 14395 7044 14399 7100
rect 14399 7044 14455 7100
rect 14455 7044 14459 7100
rect 14395 7040 14459 7044
rect 14475 7100 14539 7104
rect 14475 7044 14479 7100
rect 14479 7044 14535 7100
rect 14535 7044 14539 7100
rect 14475 7040 14539 7044
rect 14555 7100 14619 7104
rect 14555 7044 14559 7100
rect 14559 7044 14615 7100
rect 14615 7044 14619 7100
rect 14555 7040 14619 7044
rect 3521 6556 3585 6560
rect 3521 6500 3525 6556
rect 3525 6500 3581 6556
rect 3581 6500 3585 6556
rect 3521 6496 3585 6500
rect 3601 6556 3665 6560
rect 3601 6500 3605 6556
rect 3605 6500 3661 6556
rect 3661 6500 3665 6556
rect 3601 6496 3665 6500
rect 3681 6556 3745 6560
rect 3681 6500 3685 6556
rect 3685 6500 3741 6556
rect 3741 6500 3745 6556
rect 3681 6496 3745 6500
rect 3761 6556 3825 6560
rect 3761 6500 3765 6556
rect 3765 6500 3821 6556
rect 3821 6500 3825 6556
rect 3761 6496 3825 6500
rect 7339 6556 7403 6560
rect 7339 6500 7343 6556
rect 7343 6500 7399 6556
rect 7399 6500 7403 6556
rect 7339 6496 7403 6500
rect 7419 6556 7483 6560
rect 7419 6500 7423 6556
rect 7423 6500 7479 6556
rect 7479 6500 7483 6556
rect 7419 6496 7483 6500
rect 7499 6556 7563 6560
rect 7499 6500 7503 6556
rect 7503 6500 7559 6556
rect 7559 6500 7563 6556
rect 7499 6496 7563 6500
rect 7579 6556 7643 6560
rect 7579 6500 7583 6556
rect 7583 6500 7639 6556
rect 7639 6500 7643 6556
rect 7579 6496 7643 6500
rect 11157 6556 11221 6560
rect 11157 6500 11161 6556
rect 11161 6500 11217 6556
rect 11217 6500 11221 6556
rect 11157 6496 11221 6500
rect 11237 6556 11301 6560
rect 11237 6500 11241 6556
rect 11241 6500 11297 6556
rect 11297 6500 11301 6556
rect 11237 6496 11301 6500
rect 11317 6556 11381 6560
rect 11317 6500 11321 6556
rect 11321 6500 11377 6556
rect 11377 6500 11381 6556
rect 11317 6496 11381 6500
rect 11397 6556 11461 6560
rect 11397 6500 11401 6556
rect 11401 6500 11457 6556
rect 11457 6500 11461 6556
rect 11397 6496 11461 6500
rect 14975 6556 15039 6560
rect 14975 6500 14979 6556
rect 14979 6500 15035 6556
rect 15035 6500 15039 6556
rect 14975 6496 15039 6500
rect 15055 6556 15119 6560
rect 15055 6500 15059 6556
rect 15059 6500 15115 6556
rect 15115 6500 15119 6556
rect 15055 6496 15119 6500
rect 15135 6556 15199 6560
rect 15135 6500 15139 6556
rect 15139 6500 15195 6556
rect 15195 6500 15199 6556
rect 15135 6496 15199 6500
rect 15215 6556 15279 6560
rect 15215 6500 15219 6556
rect 15219 6500 15275 6556
rect 15275 6500 15279 6556
rect 15215 6496 15279 6500
rect 2861 6012 2925 6016
rect 2861 5956 2865 6012
rect 2865 5956 2921 6012
rect 2921 5956 2925 6012
rect 2861 5952 2925 5956
rect 2941 6012 3005 6016
rect 2941 5956 2945 6012
rect 2945 5956 3001 6012
rect 3001 5956 3005 6012
rect 2941 5952 3005 5956
rect 3021 6012 3085 6016
rect 3021 5956 3025 6012
rect 3025 5956 3081 6012
rect 3081 5956 3085 6012
rect 3021 5952 3085 5956
rect 3101 6012 3165 6016
rect 3101 5956 3105 6012
rect 3105 5956 3161 6012
rect 3161 5956 3165 6012
rect 3101 5952 3165 5956
rect 6679 6012 6743 6016
rect 6679 5956 6683 6012
rect 6683 5956 6739 6012
rect 6739 5956 6743 6012
rect 6679 5952 6743 5956
rect 6759 6012 6823 6016
rect 6759 5956 6763 6012
rect 6763 5956 6819 6012
rect 6819 5956 6823 6012
rect 6759 5952 6823 5956
rect 6839 6012 6903 6016
rect 6839 5956 6843 6012
rect 6843 5956 6899 6012
rect 6899 5956 6903 6012
rect 6839 5952 6903 5956
rect 6919 6012 6983 6016
rect 6919 5956 6923 6012
rect 6923 5956 6979 6012
rect 6979 5956 6983 6012
rect 6919 5952 6983 5956
rect 10497 6012 10561 6016
rect 10497 5956 10501 6012
rect 10501 5956 10557 6012
rect 10557 5956 10561 6012
rect 10497 5952 10561 5956
rect 10577 6012 10641 6016
rect 10577 5956 10581 6012
rect 10581 5956 10637 6012
rect 10637 5956 10641 6012
rect 10577 5952 10641 5956
rect 10657 6012 10721 6016
rect 10657 5956 10661 6012
rect 10661 5956 10717 6012
rect 10717 5956 10721 6012
rect 10657 5952 10721 5956
rect 10737 6012 10801 6016
rect 10737 5956 10741 6012
rect 10741 5956 10797 6012
rect 10797 5956 10801 6012
rect 10737 5952 10801 5956
rect 14315 6012 14379 6016
rect 14315 5956 14319 6012
rect 14319 5956 14375 6012
rect 14375 5956 14379 6012
rect 14315 5952 14379 5956
rect 14395 6012 14459 6016
rect 14395 5956 14399 6012
rect 14399 5956 14455 6012
rect 14455 5956 14459 6012
rect 14395 5952 14459 5956
rect 14475 6012 14539 6016
rect 14475 5956 14479 6012
rect 14479 5956 14535 6012
rect 14535 5956 14539 6012
rect 14475 5952 14539 5956
rect 14555 6012 14619 6016
rect 14555 5956 14559 6012
rect 14559 5956 14615 6012
rect 14615 5956 14619 6012
rect 14555 5952 14619 5956
rect 3521 5468 3585 5472
rect 3521 5412 3525 5468
rect 3525 5412 3581 5468
rect 3581 5412 3585 5468
rect 3521 5408 3585 5412
rect 3601 5468 3665 5472
rect 3601 5412 3605 5468
rect 3605 5412 3661 5468
rect 3661 5412 3665 5468
rect 3601 5408 3665 5412
rect 3681 5468 3745 5472
rect 3681 5412 3685 5468
rect 3685 5412 3741 5468
rect 3741 5412 3745 5468
rect 3681 5408 3745 5412
rect 3761 5468 3825 5472
rect 3761 5412 3765 5468
rect 3765 5412 3821 5468
rect 3821 5412 3825 5468
rect 3761 5408 3825 5412
rect 7339 5468 7403 5472
rect 7339 5412 7343 5468
rect 7343 5412 7399 5468
rect 7399 5412 7403 5468
rect 7339 5408 7403 5412
rect 7419 5468 7483 5472
rect 7419 5412 7423 5468
rect 7423 5412 7479 5468
rect 7479 5412 7483 5468
rect 7419 5408 7483 5412
rect 7499 5468 7563 5472
rect 7499 5412 7503 5468
rect 7503 5412 7559 5468
rect 7559 5412 7563 5468
rect 7499 5408 7563 5412
rect 7579 5468 7643 5472
rect 7579 5412 7583 5468
rect 7583 5412 7639 5468
rect 7639 5412 7643 5468
rect 7579 5408 7643 5412
rect 11157 5468 11221 5472
rect 11157 5412 11161 5468
rect 11161 5412 11217 5468
rect 11217 5412 11221 5468
rect 11157 5408 11221 5412
rect 11237 5468 11301 5472
rect 11237 5412 11241 5468
rect 11241 5412 11297 5468
rect 11297 5412 11301 5468
rect 11237 5408 11301 5412
rect 11317 5468 11381 5472
rect 11317 5412 11321 5468
rect 11321 5412 11377 5468
rect 11377 5412 11381 5468
rect 11317 5408 11381 5412
rect 11397 5468 11461 5472
rect 11397 5412 11401 5468
rect 11401 5412 11457 5468
rect 11457 5412 11461 5468
rect 11397 5408 11461 5412
rect 14975 5468 15039 5472
rect 14975 5412 14979 5468
rect 14979 5412 15035 5468
rect 15035 5412 15039 5468
rect 14975 5408 15039 5412
rect 15055 5468 15119 5472
rect 15055 5412 15059 5468
rect 15059 5412 15115 5468
rect 15115 5412 15119 5468
rect 15055 5408 15119 5412
rect 15135 5468 15199 5472
rect 15135 5412 15139 5468
rect 15139 5412 15195 5468
rect 15195 5412 15199 5468
rect 15135 5408 15199 5412
rect 15215 5468 15279 5472
rect 15215 5412 15219 5468
rect 15219 5412 15275 5468
rect 15275 5412 15279 5468
rect 15215 5408 15279 5412
rect 2861 4924 2925 4928
rect 2861 4868 2865 4924
rect 2865 4868 2921 4924
rect 2921 4868 2925 4924
rect 2861 4864 2925 4868
rect 2941 4924 3005 4928
rect 2941 4868 2945 4924
rect 2945 4868 3001 4924
rect 3001 4868 3005 4924
rect 2941 4864 3005 4868
rect 3021 4924 3085 4928
rect 3021 4868 3025 4924
rect 3025 4868 3081 4924
rect 3081 4868 3085 4924
rect 3021 4864 3085 4868
rect 3101 4924 3165 4928
rect 3101 4868 3105 4924
rect 3105 4868 3161 4924
rect 3161 4868 3165 4924
rect 3101 4864 3165 4868
rect 6679 4924 6743 4928
rect 6679 4868 6683 4924
rect 6683 4868 6739 4924
rect 6739 4868 6743 4924
rect 6679 4864 6743 4868
rect 6759 4924 6823 4928
rect 6759 4868 6763 4924
rect 6763 4868 6819 4924
rect 6819 4868 6823 4924
rect 6759 4864 6823 4868
rect 6839 4924 6903 4928
rect 6839 4868 6843 4924
rect 6843 4868 6899 4924
rect 6899 4868 6903 4924
rect 6839 4864 6903 4868
rect 6919 4924 6983 4928
rect 6919 4868 6923 4924
rect 6923 4868 6979 4924
rect 6979 4868 6983 4924
rect 6919 4864 6983 4868
rect 10497 4924 10561 4928
rect 10497 4868 10501 4924
rect 10501 4868 10557 4924
rect 10557 4868 10561 4924
rect 10497 4864 10561 4868
rect 10577 4924 10641 4928
rect 10577 4868 10581 4924
rect 10581 4868 10637 4924
rect 10637 4868 10641 4924
rect 10577 4864 10641 4868
rect 10657 4924 10721 4928
rect 10657 4868 10661 4924
rect 10661 4868 10717 4924
rect 10717 4868 10721 4924
rect 10657 4864 10721 4868
rect 10737 4924 10801 4928
rect 10737 4868 10741 4924
rect 10741 4868 10797 4924
rect 10797 4868 10801 4924
rect 10737 4864 10801 4868
rect 14315 4924 14379 4928
rect 14315 4868 14319 4924
rect 14319 4868 14375 4924
rect 14375 4868 14379 4924
rect 14315 4864 14379 4868
rect 14395 4924 14459 4928
rect 14395 4868 14399 4924
rect 14399 4868 14455 4924
rect 14455 4868 14459 4924
rect 14395 4864 14459 4868
rect 14475 4924 14539 4928
rect 14475 4868 14479 4924
rect 14479 4868 14535 4924
rect 14535 4868 14539 4924
rect 14475 4864 14539 4868
rect 14555 4924 14619 4928
rect 14555 4868 14559 4924
rect 14559 4868 14615 4924
rect 14615 4868 14619 4924
rect 14555 4864 14619 4868
rect 3521 4380 3585 4384
rect 3521 4324 3525 4380
rect 3525 4324 3581 4380
rect 3581 4324 3585 4380
rect 3521 4320 3585 4324
rect 3601 4380 3665 4384
rect 3601 4324 3605 4380
rect 3605 4324 3661 4380
rect 3661 4324 3665 4380
rect 3601 4320 3665 4324
rect 3681 4380 3745 4384
rect 3681 4324 3685 4380
rect 3685 4324 3741 4380
rect 3741 4324 3745 4380
rect 3681 4320 3745 4324
rect 3761 4380 3825 4384
rect 3761 4324 3765 4380
rect 3765 4324 3821 4380
rect 3821 4324 3825 4380
rect 3761 4320 3825 4324
rect 7339 4380 7403 4384
rect 7339 4324 7343 4380
rect 7343 4324 7399 4380
rect 7399 4324 7403 4380
rect 7339 4320 7403 4324
rect 7419 4380 7483 4384
rect 7419 4324 7423 4380
rect 7423 4324 7479 4380
rect 7479 4324 7483 4380
rect 7419 4320 7483 4324
rect 7499 4380 7563 4384
rect 7499 4324 7503 4380
rect 7503 4324 7559 4380
rect 7559 4324 7563 4380
rect 7499 4320 7563 4324
rect 7579 4380 7643 4384
rect 7579 4324 7583 4380
rect 7583 4324 7639 4380
rect 7639 4324 7643 4380
rect 7579 4320 7643 4324
rect 11157 4380 11221 4384
rect 11157 4324 11161 4380
rect 11161 4324 11217 4380
rect 11217 4324 11221 4380
rect 11157 4320 11221 4324
rect 11237 4380 11301 4384
rect 11237 4324 11241 4380
rect 11241 4324 11297 4380
rect 11297 4324 11301 4380
rect 11237 4320 11301 4324
rect 11317 4380 11381 4384
rect 11317 4324 11321 4380
rect 11321 4324 11377 4380
rect 11377 4324 11381 4380
rect 11317 4320 11381 4324
rect 11397 4380 11461 4384
rect 11397 4324 11401 4380
rect 11401 4324 11457 4380
rect 11457 4324 11461 4380
rect 11397 4320 11461 4324
rect 14975 4380 15039 4384
rect 14975 4324 14979 4380
rect 14979 4324 15035 4380
rect 15035 4324 15039 4380
rect 14975 4320 15039 4324
rect 15055 4380 15119 4384
rect 15055 4324 15059 4380
rect 15059 4324 15115 4380
rect 15115 4324 15119 4380
rect 15055 4320 15119 4324
rect 15135 4380 15199 4384
rect 15135 4324 15139 4380
rect 15139 4324 15195 4380
rect 15195 4324 15199 4380
rect 15135 4320 15199 4324
rect 15215 4380 15279 4384
rect 15215 4324 15219 4380
rect 15219 4324 15275 4380
rect 15275 4324 15279 4380
rect 15215 4320 15279 4324
rect 2861 3836 2925 3840
rect 2861 3780 2865 3836
rect 2865 3780 2921 3836
rect 2921 3780 2925 3836
rect 2861 3776 2925 3780
rect 2941 3836 3005 3840
rect 2941 3780 2945 3836
rect 2945 3780 3001 3836
rect 3001 3780 3005 3836
rect 2941 3776 3005 3780
rect 3021 3836 3085 3840
rect 3021 3780 3025 3836
rect 3025 3780 3081 3836
rect 3081 3780 3085 3836
rect 3021 3776 3085 3780
rect 3101 3836 3165 3840
rect 3101 3780 3105 3836
rect 3105 3780 3161 3836
rect 3161 3780 3165 3836
rect 3101 3776 3165 3780
rect 6679 3836 6743 3840
rect 6679 3780 6683 3836
rect 6683 3780 6739 3836
rect 6739 3780 6743 3836
rect 6679 3776 6743 3780
rect 6759 3836 6823 3840
rect 6759 3780 6763 3836
rect 6763 3780 6819 3836
rect 6819 3780 6823 3836
rect 6759 3776 6823 3780
rect 6839 3836 6903 3840
rect 6839 3780 6843 3836
rect 6843 3780 6899 3836
rect 6899 3780 6903 3836
rect 6839 3776 6903 3780
rect 6919 3836 6983 3840
rect 6919 3780 6923 3836
rect 6923 3780 6979 3836
rect 6979 3780 6983 3836
rect 6919 3776 6983 3780
rect 10497 3836 10561 3840
rect 10497 3780 10501 3836
rect 10501 3780 10557 3836
rect 10557 3780 10561 3836
rect 10497 3776 10561 3780
rect 10577 3836 10641 3840
rect 10577 3780 10581 3836
rect 10581 3780 10637 3836
rect 10637 3780 10641 3836
rect 10577 3776 10641 3780
rect 10657 3836 10721 3840
rect 10657 3780 10661 3836
rect 10661 3780 10717 3836
rect 10717 3780 10721 3836
rect 10657 3776 10721 3780
rect 10737 3836 10801 3840
rect 10737 3780 10741 3836
rect 10741 3780 10797 3836
rect 10797 3780 10801 3836
rect 10737 3776 10801 3780
rect 14315 3836 14379 3840
rect 14315 3780 14319 3836
rect 14319 3780 14375 3836
rect 14375 3780 14379 3836
rect 14315 3776 14379 3780
rect 14395 3836 14459 3840
rect 14395 3780 14399 3836
rect 14399 3780 14455 3836
rect 14455 3780 14459 3836
rect 14395 3776 14459 3780
rect 14475 3836 14539 3840
rect 14475 3780 14479 3836
rect 14479 3780 14535 3836
rect 14535 3780 14539 3836
rect 14475 3776 14539 3780
rect 14555 3836 14619 3840
rect 14555 3780 14559 3836
rect 14559 3780 14615 3836
rect 14615 3780 14619 3836
rect 14555 3776 14619 3780
rect 3521 3292 3585 3296
rect 3521 3236 3525 3292
rect 3525 3236 3581 3292
rect 3581 3236 3585 3292
rect 3521 3232 3585 3236
rect 3601 3292 3665 3296
rect 3601 3236 3605 3292
rect 3605 3236 3661 3292
rect 3661 3236 3665 3292
rect 3601 3232 3665 3236
rect 3681 3292 3745 3296
rect 3681 3236 3685 3292
rect 3685 3236 3741 3292
rect 3741 3236 3745 3292
rect 3681 3232 3745 3236
rect 3761 3292 3825 3296
rect 3761 3236 3765 3292
rect 3765 3236 3821 3292
rect 3821 3236 3825 3292
rect 3761 3232 3825 3236
rect 7339 3292 7403 3296
rect 7339 3236 7343 3292
rect 7343 3236 7399 3292
rect 7399 3236 7403 3292
rect 7339 3232 7403 3236
rect 7419 3292 7483 3296
rect 7419 3236 7423 3292
rect 7423 3236 7479 3292
rect 7479 3236 7483 3292
rect 7419 3232 7483 3236
rect 7499 3292 7563 3296
rect 7499 3236 7503 3292
rect 7503 3236 7559 3292
rect 7559 3236 7563 3292
rect 7499 3232 7563 3236
rect 7579 3292 7643 3296
rect 7579 3236 7583 3292
rect 7583 3236 7639 3292
rect 7639 3236 7643 3292
rect 7579 3232 7643 3236
rect 11157 3292 11221 3296
rect 11157 3236 11161 3292
rect 11161 3236 11217 3292
rect 11217 3236 11221 3292
rect 11157 3232 11221 3236
rect 11237 3292 11301 3296
rect 11237 3236 11241 3292
rect 11241 3236 11297 3292
rect 11297 3236 11301 3292
rect 11237 3232 11301 3236
rect 11317 3292 11381 3296
rect 11317 3236 11321 3292
rect 11321 3236 11377 3292
rect 11377 3236 11381 3292
rect 11317 3232 11381 3236
rect 11397 3292 11461 3296
rect 11397 3236 11401 3292
rect 11401 3236 11457 3292
rect 11457 3236 11461 3292
rect 11397 3232 11461 3236
rect 14975 3292 15039 3296
rect 14975 3236 14979 3292
rect 14979 3236 15035 3292
rect 15035 3236 15039 3292
rect 14975 3232 15039 3236
rect 15055 3292 15119 3296
rect 15055 3236 15059 3292
rect 15059 3236 15115 3292
rect 15115 3236 15119 3292
rect 15055 3232 15119 3236
rect 15135 3292 15199 3296
rect 15135 3236 15139 3292
rect 15139 3236 15195 3292
rect 15195 3236 15199 3292
rect 15135 3232 15199 3236
rect 15215 3292 15279 3296
rect 15215 3236 15219 3292
rect 15219 3236 15275 3292
rect 15275 3236 15279 3292
rect 15215 3232 15279 3236
rect 2861 2748 2925 2752
rect 2861 2692 2865 2748
rect 2865 2692 2921 2748
rect 2921 2692 2925 2748
rect 2861 2688 2925 2692
rect 2941 2748 3005 2752
rect 2941 2692 2945 2748
rect 2945 2692 3001 2748
rect 3001 2692 3005 2748
rect 2941 2688 3005 2692
rect 3021 2748 3085 2752
rect 3021 2692 3025 2748
rect 3025 2692 3081 2748
rect 3081 2692 3085 2748
rect 3021 2688 3085 2692
rect 3101 2748 3165 2752
rect 3101 2692 3105 2748
rect 3105 2692 3161 2748
rect 3161 2692 3165 2748
rect 3101 2688 3165 2692
rect 6679 2748 6743 2752
rect 6679 2692 6683 2748
rect 6683 2692 6739 2748
rect 6739 2692 6743 2748
rect 6679 2688 6743 2692
rect 6759 2748 6823 2752
rect 6759 2692 6763 2748
rect 6763 2692 6819 2748
rect 6819 2692 6823 2748
rect 6759 2688 6823 2692
rect 6839 2748 6903 2752
rect 6839 2692 6843 2748
rect 6843 2692 6899 2748
rect 6899 2692 6903 2748
rect 6839 2688 6903 2692
rect 6919 2748 6983 2752
rect 6919 2692 6923 2748
rect 6923 2692 6979 2748
rect 6979 2692 6983 2748
rect 6919 2688 6983 2692
rect 10497 2748 10561 2752
rect 10497 2692 10501 2748
rect 10501 2692 10557 2748
rect 10557 2692 10561 2748
rect 10497 2688 10561 2692
rect 10577 2748 10641 2752
rect 10577 2692 10581 2748
rect 10581 2692 10637 2748
rect 10637 2692 10641 2748
rect 10577 2688 10641 2692
rect 10657 2748 10721 2752
rect 10657 2692 10661 2748
rect 10661 2692 10717 2748
rect 10717 2692 10721 2748
rect 10657 2688 10721 2692
rect 10737 2748 10801 2752
rect 10737 2692 10741 2748
rect 10741 2692 10797 2748
rect 10797 2692 10801 2748
rect 10737 2688 10801 2692
rect 14315 2748 14379 2752
rect 14315 2692 14319 2748
rect 14319 2692 14375 2748
rect 14375 2692 14379 2748
rect 14315 2688 14379 2692
rect 14395 2748 14459 2752
rect 14395 2692 14399 2748
rect 14399 2692 14455 2748
rect 14455 2692 14459 2748
rect 14395 2688 14459 2692
rect 14475 2748 14539 2752
rect 14475 2692 14479 2748
rect 14479 2692 14535 2748
rect 14535 2692 14539 2748
rect 14475 2688 14539 2692
rect 14555 2748 14619 2752
rect 14555 2692 14559 2748
rect 14559 2692 14615 2748
rect 14615 2692 14619 2748
rect 14555 2688 14619 2692
rect 3521 2204 3585 2208
rect 3521 2148 3525 2204
rect 3525 2148 3581 2204
rect 3581 2148 3585 2204
rect 3521 2144 3585 2148
rect 3601 2204 3665 2208
rect 3601 2148 3605 2204
rect 3605 2148 3661 2204
rect 3661 2148 3665 2204
rect 3601 2144 3665 2148
rect 3681 2204 3745 2208
rect 3681 2148 3685 2204
rect 3685 2148 3741 2204
rect 3741 2148 3745 2204
rect 3681 2144 3745 2148
rect 3761 2204 3825 2208
rect 3761 2148 3765 2204
rect 3765 2148 3821 2204
rect 3821 2148 3825 2204
rect 3761 2144 3825 2148
rect 7339 2204 7403 2208
rect 7339 2148 7343 2204
rect 7343 2148 7399 2204
rect 7399 2148 7403 2204
rect 7339 2144 7403 2148
rect 7419 2204 7483 2208
rect 7419 2148 7423 2204
rect 7423 2148 7479 2204
rect 7479 2148 7483 2204
rect 7419 2144 7483 2148
rect 7499 2204 7563 2208
rect 7499 2148 7503 2204
rect 7503 2148 7559 2204
rect 7559 2148 7563 2204
rect 7499 2144 7563 2148
rect 7579 2204 7643 2208
rect 7579 2148 7583 2204
rect 7583 2148 7639 2204
rect 7639 2148 7643 2204
rect 7579 2144 7643 2148
rect 11157 2204 11221 2208
rect 11157 2148 11161 2204
rect 11161 2148 11217 2204
rect 11217 2148 11221 2204
rect 11157 2144 11221 2148
rect 11237 2204 11301 2208
rect 11237 2148 11241 2204
rect 11241 2148 11297 2204
rect 11297 2148 11301 2204
rect 11237 2144 11301 2148
rect 11317 2204 11381 2208
rect 11317 2148 11321 2204
rect 11321 2148 11377 2204
rect 11377 2148 11381 2204
rect 11317 2144 11381 2148
rect 11397 2204 11461 2208
rect 11397 2148 11401 2204
rect 11401 2148 11457 2204
rect 11457 2148 11461 2204
rect 11397 2144 11461 2148
rect 14975 2204 15039 2208
rect 14975 2148 14979 2204
rect 14979 2148 15035 2204
rect 15035 2148 15039 2204
rect 14975 2144 15039 2148
rect 15055 2204 15119 2208
rect 15055 2148 15059 2204
rect 15059 2148 15115 2204
rect 15115 2148 15119 2204
rect 15055 2144 15119 2148
rect 15135 2204 15199 2208
rect 15135 2148 15139 2204
rect 15139 2148 15195 2204
rect 15195 2148 15199 2204
rect 15135 2144 15199 2148
rect 15215 2204 15279 2208
rect 15215 2148 15219 2204
rect 15219 2148 15275 2204
rect 15275 2148 15279 2204
rect 15215 2144 15279 2148
<< metal4 >>
rect 2853 16896 3173 17456
rect 2853 16832 2861 16896
rect 2925 16832 2941 16896
rect 3005 16832 3021 16896
rect 3085 16832 3101 16896
rect 3165 16832 3173 16896
rect 2853 15808 3173 16832
rect 2853 15744 2861 15808
rect 2925 15744 2941 15808
rect 3005 15744 3021 15808
rect 3085 15744 3101 15808
rect 3165 15744 3173 15808
rect 2853 15622 3173 15744
rect 2853 15386 2895 15622
rect 3131 15386 3173 15622
rect 2853 14720 3173 15386
rect 2853 14656 2861 14720
rect 2925 14656 2941 14720
rect 3005 14656 3021 14720
rect 3085 14656 3101 14720
rect 3165 14656 3173 14720
rect 2853 13632 3173 14656
rect 2853 13568 2861 13632
rect 2925 13568 2941 13632
rect 3005 13568 3021 13632
rect 3085 13568 3101 13632
rect 3165 13568 3173 13632
rect 2853 12544 3173 13568
rect 2853 12480 2861 12544
rect 2925 12480 2941 12544
rect 3005 12480 3021 12544
rect 3085 12480 3101 12544
rect 3165 12480 3173 12544
rect 2853 11814 3173 12480
rect 2853 11578 2895 11814
rect 3131 11578 3173 11814
rect 2853 11456 3173 11578
rect 2853 11392 2861 11456
rect 2925 11392 2941 11456
rect 3005 11392 3021 11456
rect 3085 11392 3101 11456
rect 3165 11392 3173 11456
rect 2853 10368 3173 11392
rect 2853 10304 2861 10368
rect 2925 10304 2941 10368
rect 3005 10304 3021 10368
rect 3085 10304 3101 10368
rect 3165 10304 3173 10368
rect 2853 9280 3173 10304
rect 2853 9216 2861 9280
rect 2925 9216 2941 9280
rect 3005 9216 3021 9280
rect 3085 9216 3101 9280
rect 3165 9216 3173 9280
rect 2853 8192 3173 9216
rect 2853 8128 2861 8192
rect 2925 8128 2941 8192
rect 3005 8128 3021 8192
rect 3085 8128 3101 8192
rect 3165 8128 3173 8192
rect 2853 8006 3173 8128
rect 2853 7770 2895 8006
rect 3131 7770 3173 8006
rect 2853 7104 3173 7770
rect 2853 7040 2861 7104
rect 2925 7040 2941 7104
rect 3005 7040 3021 7104
rect 3085 7040 3101 7104
rect 3165 7040 3173 7104
rect 2853 6016 3173 7040
rect 2853 5952 2861 6016
rect 2925 5952 2941 6016
rect 3005 5952 3021 6016
rect 3085 5952 3101 6016
rect 3165 5952 3173 6016
rect 2853 4928 3173 5952
rect 2853 4864 2861 4928
rect 2925 4864 2941 4928
rect 3005 4864 3021 4928
rect 3085 4864 3101 4928
rect 3165 4864 3173 4928
rect 2853 4198 3173 4864
rect 2853 3962 2895 4198
rect 3131 3962 3173 4198
rect 2853 3840 3173 3962
rect 2853 3776 2861 3840
rect 2925 3776 2941 3840
rect 3005 3776 3021 3840
rect 3085 3776 3101 3840
rect 3165 3776 3173 3840
rect 2853 2752 3173 3776
rect 2853 2688 2861 2752
rect 2925 2688 2941 2752
rect 3005 2688 3021 2752
rect 3085 2688 3101 2752
rect 3165 2688 3173 2752
rect 2853 2128 3173 2688
rect 3513 17440 3833 17456
rect 3513 17376 3521 17440
rect 3585 17376 3601 17440
rect 3665 17376 3681 17440
rect 3745 17376 3761 17440
rect 3825 17376 3833 17440
rect 3513 16352 3833 17376
rect 3513 16288 3521 16352
rect 3585 16288 3601 16352
rect 3665 16288 3681 16352
rect 3745 16288 3761 16352
rect 3825 16288 3833 16352
rect 3513 16282 3833 16288
rect 3513 16046 3555 16282
rect 3791 16046 3833 16282
rect 3513 15264 3833 16046
rect 3513 15200 3521 15264
rect 3585 15200 3601 15264
rect 3665 15200 3681 15264
rect 3745 15200 3761 15264
rect 3825 15200 3833 15264
rect 3513 14176 3833 15200
rect 3513 14112 3521 14176
rect 3585 14112 3601 14176
rect 3665 14112 3681 14176
rect 3745 14112 3761 14176
rect 3825 14112 3833 14176
rect 3513 13088 3833 14112
rect 3513 13024 3521 13088
rect 3585 13024 3601 13088
rect 3665 13024 3681 13088
rect 3745 13024 3761 13088
rect 3825 13024 3833 13088
rect 3513 12474 3833 13024
rect 3513 12238 3555 12474
rect 3791 12238 3833 12474
rect 3513 12000 3833 12238
rect 3513 11936 3521 12000
rect 3585 11936 3601 12000
rect 3665 11936 3681 12000
rect 3745 11936 3761 12000
rect 3825 11936 3833 12000
rect 3513 10912 3833 11936
rect 3513 10848 3521 10912
rect 3585 10848 3601 10912
rect 3665 10848 3681 10912
rect 3745 10848 3761 10912
rect 3825 10848 3833 10912
rect 3513 9824 3833 10848
rect 3513 9760 3521 9824
rect 3585 9760 3601 9824
rect 3665 9760 3681 9824
rect 3745 9760 3761 9824
rect 3825 9760 3833 9824
rect 3513 8736 3833 9760
rect 3513 8672 3521 8736
rect 3585 8672 3601 8736
rect 3665 8672 3681 8736
rect 3745 8672 3761 8736
rect 3825 8672 3833 8736
rect 3513 8666 3833 8672
rect 3513 8430 3555 8666
rect 3791 8430 3833 8666
rect 3513 7648 3833 8430
rect 3513 7584 3521 7648
rect 3585 7584 3601 7648
rect 3665 7584 3681 7648
rect 3745 7584 3761 7648
rect 3825 7584 3833 7648
rect 3513 6560 3833 7584
rect 3513 6496 3521 6560
rect 3585 6496 3601 6560
rect 3665 6496 3681 6560
rect 3745 6496 3761 6560
rect 3825 6496 3833 6560
rect 3513 5472 3833 6496
rect 3513 5408 3521 5472
rect 3585 5408 3601 5472
rect 3665 5408 3681 5472
rect 3745 5408 3761 5472
rect 3825 5408 3833 5472
rect 3513 4858 3833 5408
rect 3513 4622 3555 4858
rect 3791 4622 3833 4858
rect 3513 4384 3833 4622
rect 3513 4320 3521 4384
rect 3585 4320 3601 4384
rect 3665 4320 3681 4384
rect 3745 4320 3761 4384
rect 3825 4320 3833 4384
rect 3513 3296 3833 4320
rect 3513 3232 3521 3296
rect 3585 3232 3601 3296
rect 3665 3232 3681 3296
rect 3745 3232 3761 3296
rect 3825 3232 3833 3296
rect 3513 2208 3833 3232
rect 3513 2144 3521 2208
rect 3585 2144 3601 2208
rect 3665 2144 3681 2208
rect 3745 2144 3761 2208
rect 3825 2144 3833 2208
rect 3513 2128 3833 2144
rect 6671 16896 6991 17456
rect 6671 16832 6679 16896
rect 6743 16832 6759 16896
rect 6823 16832 6839 16896
rect 6903 16832 6919 16896
rect 6983 16832 6991 16896
rect 6671 15808 6991 16832
rect 6671 15744 6679 15808
rect 6743 15744 6759 15808
rect 6823 15744 6839 15808
rect 6903 15744 6919 15808
rect 6983 15744 6991 15808
rect 6671 15622 6991 15744
rect 6671 15386 6713 15622
rect 6949 15386 6991 15622
rect 6671 14720 6991 15386
rect 6671 14656 6679 14720
rect 6743 14656 6759 14720
rect 6823 14656 6839 14720
rect 6903 14656 6919 14720
rect 6983 14656 6991 14720
rect 6671 13632 6991 14656
rect 6671 13568 6679 13632
rect 6743 13568 6759 13632
rect 6823 13568 6839 13632
rect 6903 13568 6919 13632
rect 6983 13568 6991 13632
rect 6671 12544 6991 13568
rect 6671 12480 6679 12544
rect 6743 12480 6759 12544
rect 6823 12480 6839 12544
rect 6903 12480 6919 12544
rect 6983 12480 6991 12544
rect 6671 11814 6991 12480
rect 6671 11578 6713 11814
rect 6949 11578 6991 11814
rect 6671 11456 6991 11578
rect 6671 11392 6679 11456
rect 6743 11392 6759 11456
rect 6823 11392 6839 11456
rect 6903 11392 6919 11456
rect 6983 11392 6991 11456
rect 6671 10368 6991 11392
rect 6671 10304 6679 10368
rect 6743 10304 6759 10368
rect 6823 10304 6839 10368
rect 6903 10304 6919 10368
rect 6983 10304 6991 10368
rect 6671 9280 6991 10304
rect 6671 9216 6679 9280
rect 6743 9216 6759 9280
rect 6823 9216 6839 9280
rect 6903 9216 6919 9280
rect 6983 9216 6991 9280
rect 6671 8192 6991 9216
rect 6671 8128 6679 8192
rect 6743 8128 6759 8192
rect 6823 8128 6839 8192
rect 6903 8128 6919 8192
rect 6983 8128 6991 8192
rect 6671 8006 6991 8128
rect 6671 7770 6713 8006
rect 6949 7770 6991 8006
rect 6671 7104 6991 7770
rect 6671 7040 6679 7104
rect 6743 7040 6759 7104
rect 6823 7040 6839 7104
rect 6903 7040 6919 7104
rect 6983 7040 6991 7104
rect 6671 6016 6991 7040
rect 6671 5952 6679 6016
rect 6743 5952 6759 6016
rect 6823 5952 6839 6016
rect 6903 5952 6919 6016
rect 6983 5952 6991 6016
rect 6671 4928 6991 5952
rect 6671 4864 6679 4928
rect 6743 4864 6759 4928
rect 6823 4864 6839 4928
rect 6903 4864 6919 4928
rect 6983 4864 6991 4928
rect 6671 4198 6991 4864
rect 6671 3962 6713 4198
rect 6949 3962 6991 4198
rect 6671 3840 6991 3962
rect 6671 3776 6679 3840
rect 6743 3776 6759 3840
rect 6823 3776 6839 3840
rect 6903 3776 6919 3840
rect 6983 3776 6991 3840
rect 6671 2752 6991 3776
rect 6671 2688 6679 2752
rect 6743 2688 6759 2752
rect 6823 2688 6839 2752
rect 6903 2688 6919 2752
rect 6983 2688 6991 2752
rect 6671 2128 6991 2688
rect 7331 17440 7651 17456
rect 7331 17376 7339 17440
rect 7403 17376 7419 17440
rect 7483 17376 7499 17440
rect 7563 17376 7579 17440
rect 7643 17376 7651 17440
rect 7331 16352 7651 17376
rect 7331 16288 7339 16352
rect 7403 16288 7419 16352
rect 7483 16288 7499 16352
rect 7563 16288 7579 16352
rect 7643 16288 7651 16352
rect 7331 16282 7651 16288
rect 7331 16046 7373 16282
rect 7609 16046 7651 16282
rect 7331 15264 7651 16046
rect 7331 15200 7339 15264
rect 7403 15200 7419 15264
rect 7483 15200 7499 15264
rect 7563 15200 7579 15264
rect 7643 15200 7651 15264
rect 7331 14176 7651 15200
rect 7331 14112 7339 14176
rect 7403 14112 7419 14176
rect 7483 14112 7499 14176
rect 7563 14112 7579 14176
rect 7643 14112 7651 14176
rect 7331 13088 7651 14112
rect 7331 13024 7339 13088
rect 7403 13024 7419 13088
rect 7483 13024 7499 13088
rect 7563 13024 7579 13088
rect 7643 13024 7651 13088
rect 7331 12474 7651 13024
rect 7331 12238 7373 12474
rect 7609 12238 7651 12474
rect 7331 12000 7651 12238
rect 7331 11936 7339 12000
rect 7403 11936 7419 12000
rect 7483 11936 7499 12000
rect 7563 11936 7579 12000
rect 7643 11936 7651 12000
rect 7331 10912 7651 11936
rect 7331 10848 7339 10912
rect 7403 10848 7419 10912
rect 7483 10848 7499 10912
rect 7563 10848 7579 10912
rect 7643 10848 7651 10912
rect 7331 9824 7651 10848
rect 7331 9760 7339 9824
rect 7403 9760 7419 9824
rect 7483 9760 7499 9824
rect 7563 9760 7579 9824
rect 7643 9760 7651 9824
rect 7331 8736 7651 9760
rect 7331 8672 7339 8736
rect 7403 8672 7419 8736
rect 7483 8672 7499 8736
rect 7563 8672 7579 8736
rect 7643 8672 7651 8736
rect 7331 8666 7651 8672
rect 7331 8430 7373 8666
rect 7609 8430 7651 8666
rect 7331 7648 7651 8430
rect 7331 7584 7339 7648
rect 7403 7584 7419 7648
rect 7483 7584 7499 7648
rect 7563 7584 7579 7648
rect 7643 7584 7651 7648
rect 7331 6560 7651 7584
rect 7331 6496 7339 6560
rect 7403 6496 7419 6560
rect 7483 6496 7499 6560
rect 7563 6496 7579 6560
rect 7643 6496 7651 6560
rect 7331 5472 7651 6496
rect 7331 5408 7339 5472
rect 7403 5408 7419 5472
rect 7483 5408 7499 5472
rect 7563 5408 7579 5472
rect 7643 5408 7651 5472
rect 7331 4858 7651 5408
rect 7331 4622 7373 4858
rect 7609 4622 7651 4858
rect 7331 4384 7651 4622
rect 7331 4320 7339 4384
rect 7403 4320 7419 4384
rect 7483 4320 7499 4384
rect 7563 4320 7579 4384
rect 7643 4320 7651 4384
rect 7331 3296 7651 4320
rect 7331 3232 7339 3296
rect 7403 3232 7419 3296
rect 7483 3232 7499 3296
rect 7563 3232 7579 3296
rect 7643 3232 7651 3296
rect 7331 2208 7651 3232
rect 7331 2144 7339 2208
rect 7403 2144 7419 2208
rect 7483 2144 7499 2208
rect 7563 2144 7579 2208
rect 7643 2144 7651 2208
rect 7331 2128 7651 2144
rect 10489 16896 10809 17456
rect 10489 16832 10497 16896
rect 10561 16832 10577 16896
rect 10641 16832 10657 16896
rect 10721 16832 10737 16896
rect 10801 16832 10809 16896
rect 10489 15808 10809 16832
rect 10489 15744 10497 15808
rect 10561 15744 10577 15808
rect 10641 15744 10657 15808
rect 10721 15744 10737 15808
rect 10801 15744 10809 15808
rect 10489 15622 10809 15744
rect 10489 15386 10531 15622
rect 10767 15386 10809 15622
rect 10489 14720 10809 15386
rect 10489 14656 10497 14720
rect 10561 14656 10577 14720
rect 10641 14656 10657 14720
rect 10721 14656 10737 14720
rect 10801 14656 10809 14720
rect 10489 13632 10809 14656
rect 10489 13568 10497 13632
rect 10561 13568 10577 13632
rect 10641 13568 10657 13632
rect 10721 13568 10737 13632
rect 10801 13568 10809 13632
rect 10489 12544 10809 13568
rect 10489 12480 10497 12544
rect 10561 12480 10577 12544
rect 10641 12480 10657 12544
rect 10721 12480 10737 12544
rect 10801 12480 10809 12544
rect 10489 11814 10809 12480
rect 10489 11578 10531 11814
rect 10767 11578 10809 11814
rect 10489 11456 10809 11578
rect 10489 11392 10497 11456
rect 10561 11392 10577 11456
rect 10641 11392 10657 11456
rect 10721 11392 10737 11456
rect 10801 11392 10809 11456
rect 10489 10368 10809 11392
rect 10489 10304 10497 10368
rect 10561 10304 10577 10368
rect 10641 10304 10657 10368
rect 10721 10304 10737 10368
rect 10801 10304 10809 10368
rect 10489 9280 10809 10304
rect 10489 9216 10497 9280
rect 10561 9216 10577 9280
rect 10641 9216 10657 9280
rect 10721 9216 10737 9280
rect 10801 9216 10809 9280
rect 10489 8192 10809 9216
rect 10489 8128 10497 8192
rect 10561 8128 10577 8192
rect 10641 8128 10657 8192
rect 10721 8128 10737 8192
rect 10801 8128 10809 8192
rect 10489 8006 10809 8128
rect 10489 7770 10531 8006
rect 10767 7770 10809 8006
rect 10489 7104 10809 7770
rect 10489 7040 10497 7104
rect 10561 7040 10577 7104
rect 10641 7040 10657 7104
rect 10721 7040 10737 7104
rect 10801 7040 10809 7104
rect 10489 6016 10809 7040
rect 10489 5952 10497 6016
rect 10561 5952 10577 6016
rect 10641 5952 10657 6016
rect 10721 5952 10737 6016
rect 10801 5952 10809 6016
rect 10489 4928 10809 5952
rect 10489 4864 10497 4928
rect 10561 4864 10577 4928
rect 10641 4864 10657 4928
rect 10721 4864 10737 4928
rect 10801 4864 10809 4928
rect 10489 4198 10809 4864
rect 10489 3962 10531 4198
rect 10767 3962 10809 4198
rect 10489 3840 10809 3962
rect 10489 3776 10497 3840
rect 10561 3776 10577 3840
rect 10641 3776 10657 3840
rect 10721 3776 10737 3840
rect 10801 3776 10809 3840
rect 10489 2752 10809 3776
rect 10489 2688 10497 2752
rect 10561 2688 10577 2752
rect 10641 2688 10657 2752
rect 10721 2688 10737 2752
rect 10801 2688 10809 2752
rect 10489 2128 10809 2688
rect 11149 17440 11469 17456
rect 11149 17376 11157 17440
rect 11221 17376 11237 17440
rect 11301 17376 11317 17440
rect 11381 17376 11397 17440
rect 11461 17376 11469 17440
rect 11149 16352 11469 17376
rect 11149 16288 11157 16352
rect 11221 16288 11237 16352
rect 11301 16288 11317 16352
rect 11381 16288 11397 16352
rect 11461 16288 11469 16352
rect 11149 16282 11469 16288
rect 11149 16046 11191 16282
rect 11427 16046 11469 16282
rect 11149 15264 11469 16046
rect 11149 15200 11157 15264
rect 11221 15200 11237 15264
rect 11301 15200 11317 15264
rect 11381 15200 11397 15264
rect 11461 15200 11469 15264
rect 11149 14176 11469 15200
rect 11149 14112 11157 14176
rect 11221 14112 11237 14176
rect 11301 14112 11317 14176
rect 11381 14112 11397 14176
rect 11461 14112 11469 14176
rect 11149 13088 11469 14112
rect 11149 13024 11157 13088
rect 11221 13024 11237 13088
rect 11301 13024 11317 13088
rect 11381 13024 11397 13088
rect 11461 13024 11469 13088
rect 11149 12474 11469 13024
rect 11149 12238 11191 12474
rect 11427 12238 11469 12474
rect 11149 12000 11469 12238
rect 11149 11936 11157 12000
rect 11221 11936 11237 12000
rect 11301 11936 11317 12000
rect 11381 11936 11397 12000
rect 11461 11936 11469 12000
rect 11149 10912 11469 11936
rect 11149 10848 11157 10912
rect 11221 10848 11237 10912
rect 11301 10848 11317 10912
rect 11381 10848 11397 10912
rect 11461 10848 11469 10912
rect 11149 9824 11469 10848
rect 11149 9760 11157 9824
rect 11221 9760 11237 9824
rect 11301 9760 11317 9824
rect 11381 9760 11397 9824
rect 11461 9760 11469 9824
rect 11149 8736 11469 9760
rect 11149 8672 11157 8736
rect 11221 8672 11237 8736
rect 11301 8672 11317 8736
rect 11381 8672 11397 8736
rect 11461 8672 11469 8736
rect 11149 8666 11469 8672
rect 11149 8430 11191 8666
rect 11427 8430 11469 8666
rect 11149 7648 11469 8430
rect 11149 7584 11157 7648
rect 11221 7584 11237 7648
rect 11301 7584 11317 7648
rect 11381 7584 11397 7648
rect 11461 7584 11469 7648
rect 11149 6560 11469 7584
rect 11149 6496 11157 6560
rect 11221 6496 11237 6560
rect 11301 6496 11317 6560
rect 11381 6496 11397 6560
rect 11461 6496 11469 6560
rect 11149 5472 11469 6496
rect 11149 5408 11157 5472
rect 11221 5408 11237 5472
rect 11301 5408 11317 5472
rect 11381 5408 11397 5472
rect 11461 5408 11469 5472
rect 11149 4858 11469 5408
rect 11149 4622 11191 4858
rect 11427 4622 11469 4858
rect 11149 4384 11469 4622
rect 11149 4320 11157 4384
rect 11221 4320 11237 4384
rect 11301 4320 11317 4384
rect 11381 4320 11397 4384
rect 11461 4320 11469 4384
rect 11149 3296 11469 4320
rect 11149 3232 11157 3296
rect 11221 3232 11237 3296
rect 11301 3232 11317 3296
rect 11381 3232 11397 3296
rect 11461 3232 11469 3296
rect 11149 2208 11469 3232
rect 11149 2144 11157 2208
rect 11221 2144 11237 2208
rect 11301 2144 11317 2208
rect 11381 2144 11397 2208
rect 11461 2144 11469 2208
rect 11149 2128 11469 2144
rect 14307 16896 14627 17456
rect 14307 16832 14315 16896
rect 14379 16832 14395 16896
rect 14459 16832 14475 16896
rect 14539 16832 14555 16896
rect 14619 16832 14627 16896
rect 14307 15808 14627 16832
rect 14307 15744 14315 15808
rect 14379 15744 14395 15808
rect 14459 15744 14475 15808
rect 14539 15744 14555 15808
rect 14619 15744 14627 15808
rect 14307 15622 14627 15744
rect 14307 15386 14349 15622
rect 14585 15386 14627 15622
rect 14307 14720 14627 15386
rect 14307 14656 14315 14720
rect 14379 14656 14395 14720
rect 14459 14656 14475 14720
rect 14539 14656 14555 14720
rect 14619 14656 14627 14720
rect 14307 13632 14627 14656
rect 14307 13568 14315 13632
rect 14379 13568 14395 13632
rect 14459 13568 14475 13632
rect 14539 13568 14555 13632
rect 14619 13568 14627 13632
rect 14307 12544 14627 13568
rect 14307 12480 14315 12544
rect 14379 12480 14395 12544
rect 14459 12480 14475 12544
rect 14539 12480 14555 12544
rect 14619 12480 14627 12544
rect 14307 11814 14627 12480
rect 14307 11578 14349 11814
rect 14585 11578 14627 11814
rect 14307 11456 14627 11578
rect 14307 11392 14315 11456
rect 14379 11392 14395 11456
rect 14459 11392 14475 11456
rect 14539 11392 14555 11456
rect 14619 11392 14627 11456
rect 14307 10368 14627 11392
rect 14307 10304 14315 10368
rect 14379 10304 14395 10368
rect 14459 10304 14475 10368
rect 14539 10304 14555 10368
rect 14619 10304 14627 10368
rect 14307 9280 14627 10304
rect 14307 9216 14315 9280
rect 14379 9216 14395 9280
rect 14459 9216 14475 9280
rect 14539 9216 14555 9280
rect 14619 9216 14627 9280
rect 14307 8192 14627 9216
rect 14307 8128 14315 8192
rect 14379 8128 14395 8192
rect 14459 8128 14475 8192
rect 14539 8128 14555 8192
rect 14619 8128 14627 8192
rect 14307 8006 14627 8128
rect 14307 7770 14349 8006
rect 14585 7770 14627 8006
rect 14307 7104 14627 7770
rect 14307 7040 14315 7104
rect 14379 7040 14395 7104
rect 14459 7040 14475 7104
rect 14539 7040 14555 7104
rect 14619 7040 14627 7104
rect 14307 6016 14627 7040
rect 14307 5952 14315 6016
rect 14379 5952 14395 6016
rect 14459 5952 14475 6016
rect 14539 5952 14555 6016
rect 14619 5952 14627 6016
rect 14307 4928 14627 5952
rect 14307 4864 14315 4928
rect 14379 4864 14395 4928
rect 14459 4864 14475 4928
rect 14539 4864 14555 4928
rect 14619 4864 14627 4928
rect 14307 4198 14627 4864
rect 14307 3962 14349 4198
rect 14585 3962 14627 4198
rect 14307 3840 14627 3962
rect 14307 3776 14315 3840
rect 14379 3776 14395 3840
rect 14459 3776 14475 3840
rect 14539 3776 14555 3840
rect 14619 3776 14627 3840
rect 14307 2752 14627 3776
rect 14307 2688 14315 2752
rect 14379 2688 14395 2752
rect 14459 2688 14475 2752
rect 14539 2688 14555 2752
rect 14619 2688 14627 2752
rect 14307 2128 14627 2688
rect 14967 17440 15287 17456
rect 14967 17376 14975 17440
rect 15039 17376 15055 17440
rect 15119 17376 15135 17440
rect 15199 17376 15215 17440
rect 15279 17376 15287 17440
rect 14967 16352 15287 17376
rect 14967 16288 14975 16352
rect 15039 16288 15055 16352
rect 15119 16288 15135 16352
rect 15199 16288 15215 16352
rect 15279 16288 15287 16352
rect 14967 16282 15287 16288
rect 14967 16046 15009 16282
rect 15245 16046 15287 16282
rect 14967 15264 15287 16046
rect 14967 15200 14975 15264
rect 15039 15200 15055 15264
rect 15119 15200 15135 15264
rect 15199 15200 15215 15264
rect 15279 15200 15287 15264
rect 14967 14176 15287 15200
rect 14967 14112 14975 14176
rect 15039 14112 15055 14176
rect 15119 14112 15135 14176
rect 15199 14112 15215 14176
rect 15279 14112 15287 14176
rect 14967 13088 15287 14112
rect 14967 13024 14975 13088
rect 15039 13024 15055 13088
rect 15119 13024 15135 13088
rect 15199 13024 15215 13088
rect 15279 13024 15287 13088
rect 14967 12474 15287 13024
rect 14967 12238 15009 12474
rect 15245 12238 15287 12474
rect 14967 12000 15287 12238
rect 14967 11936 14975 12000
rect 15039 11936 15055 12000
rect 15119 11936 15135 12000
rect 15199 11936 15215 12000
rect 15279 11936 15287 12000
rect 14967 10912 15287 11936
rect 14967 10848 14975 10912
rect 15039 10848 15055 10912
rect 15119 10848 15135 10912
rect 15199 10848 15215 10912
rect 15279 10848 15287 10912
rect 14967 9824 15287 10848
rect 14967 9760 14975 9824
rect 15039 9760 15055 9824
rect 15119 9760 15135 9824
rect 15199 9760 15215 9824
rect 15279 9760 15287 9824
rect 14967 8736 15287 9760
rect 14967 8672 14975 8736
rect 15039 8672 15055 8736
rect 15119 8672 15135 8736
rect 15199 8672 15215 8736
rect 15279 8672 15287 8736
rect 14967 8666 15287 8672
rect 14967 8430 15009 8666
rect 15245 8430 15287 8666
rect 14967 7648 15287 8430
rect 14967 7584 14975 7648
rect 15039 7584 15055 7648
rect 15119 7584 15135 7648
rect 15199 7584 15215 7648
rect 15279 7584 15287 7648
rect 14967 6560 15287 7584
rect 14967 6496 14975 6560
rect 15039 6496 15055 6560
rect 15119 6496 15135 6560
rect 15199 6496 15215 6560
rect 15279 6496 15287 6560
rect 14967 5472 15287 6496
rect 14967 5408 14975 5472
rect 15039 5408 15055 5472
rect 15119 5408 15135 5472
rect 15199 5408 15215 5472
rect 15279 5408 15287 5472
rect 14967 4858 15287 5408
rect 14967 4622 15009 4858
rect 15245 4622 15287 4858
rect 14967 4384 15287 4622
rect 14967 4320 14975 4384
rect 15039 4320 15055 4384
rect 15119 4320 15135 4384
rect 15199 4320 15215 4384
rect 15279 4320 15287 4384
rect 14967 3296 15287 4320
rect 14967 3232 14975 3296
rect 15039 3232 15055 3296
rect 15119 3232 15135 3296
rect 15199 3232 15215 3296
rect 15279 3232 15287 3296
rect 14967 2208 15287 3232
rect 14967 2144 14975 2208
rect 15039 2144 15055 2208
rect 15119 2144 15135 2208
rect 15199 2144 15215 2208
rect 15279 2144 15287 2208
rect 14967 2128 15287 2144
<< via4 >>
rect 2895 15386 3131 15622
rect 2895 11578 3131 11814
rect 2895 7770 3131 8006
rect 2895 3962 3131 4198
rect 3555 16046 3791 16282
rect 3555 12238 3791 12474
rect 3555 8430 3791 8666
rect 3555 4622 3791 4858
rect 6713 15386 6949 15622
rect 6713 11578 6949 11814
rect 6713 7770 6949 8006
rect 6713 3962 6949 4198
rect 7373 16046 7609 16282
rect 7373 12238 7609 12474
rect 7373 8430 7609 8666
rect 7373 4622 7609 4858
rect 10531 15386 10767 15622
rect 10531 11578 10767 11814
rect 10531 7770 10767 8006
rect 10531 3962 10767 4198
rect 11191 16046 11427 16282
rect 11191 12238 11427 12474
rect 11191 8430 11427 8666
rect 11191 4622 11427 4858
rect 14349 15386 14585 15622
rect 14349 11578 14585 11814
rect 14349 7770 14585 8006
rect 14349 3962 14585 4198
rect 15009 16046 15245 16282
rect 15009 12238 15245 12474
rect 15009 8430 15245 8666
rect 15009 4622 15245 4858
<< metal5 >>
rect 1056 16282 16424 16324
rect 1056 16046 3555 16282
rect 3791 16046 7373 16282
rect 7609 16046 11191 16282
rect 11427 16046 15009 16282
rect 15245 16046 16424 16282
rect 1056 16004 16424 16046
rect 1056 15622 16424 15664
rect 1056 15386 2895 15622
rect 3131 15386 6713 15622
rect 6949 15386 10531 15622
rect 10767 15386 14349 15622
rect 14585 15386 16424 15622
rect 1056 15344 16424 15386
rect 1056 12474 16424 12516
rect 1056 12238 3555 12474
rect 3791 12238 7373 12474
rect 7609 12238 11191 12474
rect 11427 12238 15009 12474
rect 15245 12238 16424 12474
rect 1056 12196 16424 12238
rect 1056 11814 16424 11856
rect 1056 11578 2895 11814
rect 3131 11578 6713 11814
rect 6949 11578 10531 11814
rect 10767 11578 14349 11814
rect 14585 11578 16424 11814
rect 1056 11536 16424 11578
rect 1056 8666 16424 8708
rect 1056 8430 3555 8666
rect 3791 8430 7373 8666
rect 7609 8430 11191 8666
rect 11427 8430 15009 8666
rect 15245 8430 16424 8666
rect 1056 8388 16424 8430
rect 1056 8006 16424 8048
rect 1056 7770 2895 8006
rect 3131 7770 6713 8006
rect 6949 7770 10531 8006
rect 10767 7770 14349 8006
rect 14585 7770 16424 8006
rect 1056 7728 16424 7770
rect 1056 4858 16424 4900
rect 1056 4622 3555 4858
rect 3791 4622 7373 4858
rect 7609 4622 11191 4858
rect 11427 4622 15009 4858
rect 15245 4622 16424 4858
rect 1056 4580 16424 4622
rect 1056 4198 16424 4240
rect 1056 3962 2895 4198
rect 3131 3962 6713 4198
rect 6949 3962 10531 4198
rect 10767 3962 14349 4198
rect 14585 3962 16424 4198
rect 1056 3920 16424 3962
use sky130_fd_sc_hd__xor2_1  _314_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 2300 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _315_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _316_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 6440 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _317_
timestamp 1694700623
transform -1 0 5888 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _318_
timestamp 1694700623
transform 1 0 3220 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _319_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3220 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _320_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3496 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _321_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 5060 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _322_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3680 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _323_
timestamp 1694700623
transform 1 0 4508 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _324_
timestamp 1694700623
transform 1 0 7268 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _325_
timestamp 1694700623
transform 1 0 10580 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _326_
timestamp 1694700623
transform 1 0 11040 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _327_
timestamp 1694700623
transform 1 0 11868 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _328_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 13064 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _329_
timestamp 1694700623
transform 1 0 10948 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _330_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 11776 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _331_
timestamp 1694700623
transform 1 0 12052 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _332_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 7544 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _333_
timestamp 1694700623
transform 1 0 7360 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _334_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 8832 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _335_
timestamp 1694700623
transform 1 0 8924 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _336_
timestamp 1694700623
transform 1 0 7912 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _337_
timestamp 1694700623
transform 1 0 9200 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _338_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 10212 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _339_
timestamp 1694700623
transform -1 0 11684 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _340_
timestamp 1694700623
transform 1 0 11500 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _341_
timestamp 1694700623
transform 1 0 12052 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _342_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 12420 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _343_
timestamp 1694700623
transform 1 0 12236 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _344_
timestamp 1694700623
transform -1 0 12972 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _345_
timestamp 1694700623
transform 1 0 13156 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _346_
timestamp 1694700623
transform 1 0 14260 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _347_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 14444 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _348_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 15456 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _349_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 7544 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1694700623
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _351_
timestamp 1694700623
transform 1 0 8280 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _352_
timestamp 1694700623
transform 1 0 9568 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _353_
timestamp 1694700623
transform 1 0 5520 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _354_
timestamp 1694700623
transform 1 0 2484 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _355_
timestamp 1694700623
transform 1 0 2944 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _356_
timestamp 1694700623
transform 1 0 3220 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _357_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 2760 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _358_
timestamp 1694700623
transform -1 0 4876 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _359_
timestamp 1694700623
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _360_
timestamp 1694700623
transform 1 0 4140 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _361_
timestamp 1694700623
transform 1 0 4876 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _362_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5796 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _363_
timestamp 1694700623
transform -1 0 4876 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _364_
timestamp 1694700623
transform -1 0 4508 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _365_
timestamp 1694700623
transform -1 0 4416 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _366_
timestamp 1694700623
transform 1 0 4508 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _367_
timestamp 1694700623
transform 1 0 9844 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _368_
timestamp 1694700623
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _369_
timestamp 1694700623
transform 1 0 11408 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _370_
timestamp 1694700623
transform 1 0 12144 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _371_
timestamp 1694700623
transform 1 0 13156 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _372_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 9660 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _373_
timestamp 1694700623
transform 1 0 7084 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _374_
timestamp 1694700623
transform 1 0 7728 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _375_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 8556 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _376_
timestamp 1694700623
transform 1 0 8096 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _377_
timestamp 1694700623
transform -1 0 8556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _378_
timestamp 1694700623
transform 1 0 10396 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _379_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 10856 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _380_
timestamp 1694700623
transform 1 0 11500 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _381_
timestamp 1694700623
transform 1 0 11960 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _382_
timestamp 1694700623
transform 1 0 12328 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _383_
timestamp 1694700623
transform 1 0 12788 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _384_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 13432 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _385_
timestamp 1694700623
transform 1 0 14628 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _386_
timestamp 1694700623
transform -1 0 14904 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _387_
timestamp 1694700623
transform 1 0 14904 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _388_
timestamp 1694700623
transform 1 0 10488 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _389_
timestamp 1694700623
transform 1 0 7636 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _390_
timestamp 1694700623
transform 1 0 8372 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _391_
timestamp 1694700623
transform 1 0 8924 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _392_
timestamp 1694700623
transform 1 0 7452 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _393_
timestamp 1694700623
transform 1 0 10120 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _394_
timestamp 1694700623
transform 1 0 10120 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _395_
timestamp 1694700623
transform 1 0 10672 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _396_
timestamp 1694700623
transform 1 0 3772 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _397_
timestamp 1694700623
transform -1 0 4324 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _398_
timestamp 1694700623
transform -1 0 4784 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _399_
timestamp 1694700623
transform -1 0 5428 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _400_
timestamp 1694700623
transform 1 0 4968 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _401_
timestamp 1694700623
transform 1 0 5888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _402_
timestamp 1694700623
transform 1 0 11500 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _403_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 12420 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _404_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 12420 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _405_
timestamp 1694700623
transform 1 0 12788 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _406_
timestamp 1694700623
transform 1 0 12972 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _407_
timestamp 1694700623
transform 1 0 9016 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _408_
timestamp 1694700623
transform 1 0 10212 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _409_
timestamp 1694700623
transform -1 0 9660 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _410_
timestamp 1694700623
transform -1 0 12420 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _411_
timestamp 1694700623
transform 1 0 12420 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _412_
timestamp 1694700623
transform 1 0 12512 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _413_
timestamp 1694700623
transform 1 0 13156 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _414_
timestamp 1694700623
transform 1 0 14168 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _415_
timestamp 1694700623
transform 1 0 15088 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _416_
timestamp 1694700623
transform 1 0 14352 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _417_
timestamp 1694700623
transform 1 0 14812 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _418_
timestamp 1694700623
transform -1 0 11684 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _419_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 7360 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _420_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 7360 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _421_
timestamp 1694700623
transform 1 0 7176 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _422_
timestamp 1694700623
transform 1 0 7728 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _423_
timestamp 1694700623
transform 1 0 7912 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _424_
timestamp 1694700623
transform -1 0 7728 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _425_
timestamp 1694700623
transform 1 0 8188 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _426_
timestamp 1694700623
transform -1 0 9292 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _427_
timestamp 1694700623
transform 1 0 9016 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _428_
timestamp 1694700623
transform 1 0 9476 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _429_
timestamp 1694700623
transform 1 0 10580 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _430_
timestamp 1694700623
transform 1 0 10672 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _431_
timestamp 1694700623
transform 1 0 11040 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _432_
timestamp 1694700623
transform 1 0 5428 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _433_
timestamp 1694700623
transform 1 0 11684 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _434_
timestamp 1694700623
transform 1 0 12144 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _435_
timestamp 1694700623
transform 1 0 12788 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _436_
timestamp 1694700623
transform 1 0 13248 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _437_
timestamp 1694700623
transform -1 0 13708 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _438_
timestamp 1694700623
transform 1 0 9660 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _439_
timestamp 1694700623
transform 1 0 12972 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _440_
timestamp 1694700623
transform 1 0 13248 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _441_
timestamp 1694700623
transform 1 0 14352 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _442_
timestamp 1694700623
transform 1 0 13432 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _443_
timestamp 1694700623
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _444_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 12328 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _445_
timestamp 1694700623
transform 1 0 9660 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _446_
timestamp 1694700623
transform 1 0 7268 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _447_
timestamp 1694700623
transform -1 0 7452 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _448_
timestamp 1694700623
transform 1 0 7544 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _449_
timestamp 1694700623
transform 1 0 8372 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _450_
timestamp 1694700623
transform 1 0 8924 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _451_
timestamp 1694700623
transform -1 0 9844 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _452_
timestamp 1694700623
transform 1 0 9108 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _453_
timestamp 1694700623
transform 1 0 9844 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _454_
timestamp 1694700623
transform 1 0 10120 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _455_
timestamp 1694700623
transform 1 0 10488 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _456_
timestamp 1694700623
transform 1 0 10948 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _457_
timestamp 1694700623
transform -1 0 13064 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _458_
timestamp 1694700623
transform 1 0 13064 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _459_
timestamp 1694700623
transform -1 0 14444 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _460_
timestamp 1694700623
transform 1 0 13524 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _461_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 8280 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _462_
timestamp 1694700623
transform -1 0 6992 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _463_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5612 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _464_
timestamp 1694700623
transform 1 0 6716 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _465_
timestamp 1694700623
transform 1 0 6532 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _466_
timestamp 1694700623
transform -1 0 6716 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _467_
timestamp 1694700623
transform 1 0 7176 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _468_
timestamp 1694700623
transform 1 0 8924 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _469_
timestamp 1694700623
transform 1 0 10028 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _470_
timestamp 1694700623
transform 1 0 10212 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _471_
timestamp 1694700623
transform 1 0 11132 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _472_
timestamp 1694700623
transform -1 0 14444 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _473_
timestamp 1694700623
transform 1 0 14076 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _474_
timestamp 1694700623
transform -1 0 14076 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _475_
timestamp 1694700623
transform 1 0 9568 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _476_
timestamp 1694700623
transform 1 0 7268 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _477_
timestamp 1694700623
transform 1 0 8280 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _478_
timestamp 1694700623
transform -1 0 8280 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _479_
timestamp 1694700623
transform -1 0 10672 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _480_
timestamp 1694700623
transform 1 0 10672 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _481_
timestamp 1694700623
transform 1 0 11500 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _482_
timestamp 1694700623
transform 1 0 11684 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _483_
timestamp 1694700623
transform 1 0 12604 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _484_
timestamp 1694700623
transform 1 0 12880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _485_
timestamp 1694700623
transform 1 0 12788 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _486_
timestamp 1694700623
transform 1 0 6900 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _487_
timestamp 1694700623
transform 1 0 12144 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _488_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 12144 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _489_
timestamp 1694700623
transform 1 0 11500 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _490_
timestamp 1694700623
transform 1 0 14076 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _491_
timestamp 1694700623
transform 1 0 14720 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _492_
timestamp 1694700623
transform 1 0 15088 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _493_
timestamp 1694700623
transform 1 0 15272 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _494_
timestamp 1694700623
transform -1 0 7636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _495_
timestamp 1694700623
transform 1 0 8556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _496_
timestamp 1694700623
transform 1 0 2944 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _497_
timestamp 1694700623
transform 1 0 3496 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _498_
timestamp 1694700623
transform 1 0 2944 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _499_
timestamp 1694700623
transform -1 0 1840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _500_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1748 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _501_
timestamp 1694700623
transform -1 0 2668 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _502_
timestamp 1694700623
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _503_
timestamp 1694700623
transform 1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _504_
timestamp 1694700623
transform -1 0 2392 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _505_
timestamp 1694700623
transform 1 0 1748 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _506_
timestamp 1694700623
transform -1 0 2392 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  _507_
timestamp 1694700623
transform 1 0 2760 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _508_
timestamp 1694700623
transform -1 0 3956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_4  _509_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 2668 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _510_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 2576 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _511_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3680 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _512_
timestamp 1694700623
transform 1 0 3956 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _513_
timestamp 1694700623
transform -1 0 3680 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _514_
timestamp 1694700623
transform 1 0 2852 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _515_
timestamp 1694700623
transform 1 0 4416 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _516_
timestamp 1694700623
transform 1 0 7268 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _517_
timestamp 1694700623
transform 1 0 8004 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _518_
timestamp 1694700623
transform -1 0 4140 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _519_
timestamp 1694700623
transform -1 0 4968 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _520_
timestamp 1694700623
transform -1 0 4692 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _521_
timestamp 1694700623
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _522_
timestamp 1694700623
transform -1 0 5980 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _523_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 2392 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_2  _524_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 3128 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _525_
timestamp 1694700623
transform 1 0 1564 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _526_
timestamp 1694700623
transform 1 0 1932 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _527_
timestamp 1694700623
transform -1 0 2760 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _528_
timestamp 1694700623
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _529_
timestamp 1694700623
transform 1 0 2576 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _530_
timestamp 1694700623
transform 1 0 3220 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _531_
timestamp 1694700623
transform -1 0 4692 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _532_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 4968 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _533_
timestamp 1694700623
transform 1 0 4968 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _534_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 4324 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _535_
timestamp 1694700623
transform 1 0 2760 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _536_
timestamp 1694700623
transform -1 0 4876 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _537_
timestamp 1694700623
transform 1 0 3956 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _538_
timestamp 1694700623
transform 1 0 4968 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _539_
timestamp 1694700623
transform 1 0 5612 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _540_
timestamp 1694700623
transform 1 0 8096 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _541_
timestamp 1694700623
transform -1 0 7268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _542_
timestamp 1694700623
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _543_
timestamp 1694700623
transform 1 0 7636 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _544_
timestamp 1694700623
transform 1 0 12144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _545_
timestamp 1694700623
transform -1 0 6256 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _546_
timestamp 1694700623
transform -1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _547_
timestamp 1694700623
transform 1 0 5888 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _548_
timestamp 1694700623
transform 1 0 6532 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _549_
timestamp 1694700623
transform 1 0 8832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _550_
timestamp 1694700623
transform 1 0 7084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _551_
timestamp 1694700623
transform -1 0 9476 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _552_
timestamp 1694700623
transform -1 0 9292 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _553_
timestamp 1694700623
transform 1 0 7636 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _554_
timestamp 1694700623
transform -1 0 9200 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _555_
timestamp 1694700623
transform -1 0 6716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _556_
timestamp 1694700623
transform 1 0 6716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _557_
timestamp 1694700623
transform -1 0 6440 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _558_
timestamp 1694700623
transform 1 0 3772 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _559_
timestamp 1694700623
transform 1 0 3220 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _560_
timestamp 1694700623
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _561_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 6072 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _562_
timestamp 1694700623
transform -1 0 5888 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _563_
timestamp 1694700623
transform -1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _564_
timestamp 1694700623
transform 1 0 4784 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _565_
timestamp 1694700623
transform 1 0 6808 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _566_
timestamp 1694700623
transform 1 0 6164 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _567_
timestamp 1694700623
transform -1 0 6164 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _568_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 7728 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _569_
timestamp 1694700623
transform 1 0 7176 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _570_
timestamp 1694700623
transform 1 0 8556 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _571_
timestamp 1694700623
transform 1 0 9200 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _572_
timestamp 1694700623
transform 1 0 10028 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _573_
timestamp 1694700623
transform -1 0 10580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _574_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _575_
timestamp 1694700623
transform -1 0 2484 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _576_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5888 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _577_
timestamp 1694700623
transform -1 0 5704 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _578_
timestamp 1694700623
transform -1 0 5244 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _579_
timestamp 1694700623
transform -1 0 3312 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _580_
timestamp 1694700623
transform -1 0 4416 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _581_
timestamp 1694700623
transform 1 0 3496 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _582_
timestamp 1694700623
transform 1 0 9200 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _583_
timestamp 1694700623
transform 1 0 9292 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _584_
timestamp 1694700623
transform -1 0 7084 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _585_
timestamp 1694700623
transform 1 0 8924 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _586_
timestamp 1694700623
transform 1 0 9384 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _587_
timestamp 1694700623
transform 1 0 7912 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _588_
timestamp 1694700623
transform 1 0 8188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _589_
timestamp 1694700623
transform 1 0 10672 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _590_
timestamp 1694700623
transform -1 0 10672 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _591_
timestamp 1694700623
transform 1 0 11500 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _592_
timestamp 1694700623
transform 1 0 6992 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _593_
timestamp 1694700623
transform 1 0 6532 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _594_
timestamp 1694700623
transform -1 0 6440 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _595_
timestamp 1694700623
transform 1 0 9936 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _596_
timestamp 1694700623
transform 1 0 10304 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _597_
timestamp 1694700623
transform 1 0 11776 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _598_
timestamp 1694700623
transform 1 0 12512 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _599_
timestamp 1694700623
transform 1 0 13340 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _600_
timestamp 1694700623
transform 1 0 13524 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _601_
timestamp 1694700623
transform -1 0 14536 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _602_
timestamp 1694700623
transform -1 0 2760 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _603_
timestamp 1694700623
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_1  _604_
timestamp 1694700623
transform -1 0 1932 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _605_
timestamp 1694700623
transform -1 0 2484 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _606_
timestamp 1694700623
transform -1 0 5704 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _607_
timestamp 1694700623
transform 1 0 6992 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _608_
timestamp 1694700623
transform -1 0 6992 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _609_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5612 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _610_
timestamp 1694700623
transform 1 0 5152 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _611_
timestamp 1694700623
transform -1 0 5152 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _612_
timestamp 1694700623
transform 1 0 5152 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _613_
timestamp 1694700623
transform 1 0 1840 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _614_
timestamp 1694700623
transform -1 0 3496 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _615_
timestamp 1694700623
transform 1 0 3772 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _616_
timestamp 1694700623
transform 1 0 4232 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _617_
timestamp 1694700623
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _618_
timestamp 1694700623
transform -1 0 12972 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _619_
timestamp 1694700623
transform 1 0 6348 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _620_
timestamp 1694700623
transform 1 0 10948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _621_
timestamp 1694700623
transform 1 0 7268 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _622_
timestamp 1694700623
transform -1 0 8924 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _623_
timestamp 1694700623
transform 1 0 8832 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _624_
timestamp 1694700623
transform 1 0 7084 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _625_
timestamp 1694700623
transform 1 0 9752 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _626_
timestamp 1694700623
transform 1 0 8280 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _627_
timestamp 1694700623
transform 1 0 8924 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _628_
timestamp 1694700623
transform -1 0 8832 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _629_
timestamp 1694700623
transform 1 0 9476 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _630_
timestamp 1694700623
transform 1 0 9292 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _631_
timestamp 1694700623
transform 1 0 10120 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _632_
timestamp 1694700623
transform 1 0 10580 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _633_
timestamp 1694700623
transform 1 0 11500 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _634_
timestamp 1694700623
transform -1 0 11960 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _635_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 11960 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_4  _636_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 12788 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _637_
timestamp 1694700623
transform 1 0 12788 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _638_
timestamp 1694700623
transform 1 0 14076 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _639_
timestamp 1694700623
transform 1 0 13892 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _640_
timestamp 1694700623
transform -1 0 14904 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _641_
timestamp 1694700623
transform 1 0 2484 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _642_
timestamp 1694700623
transform 1 0 2484 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _643_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1656 0 1 11968
box -38 -48 682 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1694700623
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_37
timestamp 1694700623
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_44
timestamp 1694700623
transform 1 0 5152 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_57
timestamp 1694700623
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_65
timestamp 1694700623
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_69 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_90
timestamp 1694700623
transform 1 0 9384 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_98
timestamp 1694700623
transform 1 0 10120 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_103
timestamp 1694700623
transform 1 0 10580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1694700623
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_113
timestamp 1694700623
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_121
timestamp 1694700623
transform 1 0 12236 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_128
timestamp 1694700623
transform 1 0 12880 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1694700623
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_153
timestamp 1694700623
transform 1 0 15180 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_161
timestamp 1694700623
transform 1 0 15916 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_19
timestamp 1694700623
transform 1 0 2852 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_39
timestamp 1694700623
transform 1 0 4692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_87
timestamp 1694700623
transform 1 0 9108 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_95
timestamp 1694700623
transform 1 0 9844 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_104
timestamp 1694700623
transform 1 0 10672 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_123
timestamp 1694700623
transform 1 0 12420 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_135
timestamp 1694700623
transform 1 0 13524 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_147
timestamp 1694700623
transform 1 0 14628 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_159
timestamp 1694700623
transform 1 0 15732 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_9
timestamp 1694700623
transform 1 0 1932 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_21
timestamp 1694700623
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1694700623
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_29
timestamp 1694700623
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_36
timestamp 1694700623
transform 1 0 4416 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_48
timestamp 1694700623
transform 1 0 5520 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_64
timestamp 1694700623
transform 1 0 6992 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_72
timestamp 1694700623
transform 1 0 7728 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1694700623
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1694700623
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_85
timestamp 1694700623
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_93
timestamp 1694700623
transform 1 0 9660 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_105
timestamp 1694700623
transform 1 0 10764 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_117
timestamp 1694700623
transform 1 0 11868 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_123
timestamp 1694700623
transform 1 0 12420 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_131
timestamp 1694700623
transform 1 0 13156 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_148
timestamp 1694700623
transform 1 0 14720 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_156
timestamp 1694700623
transform 1 0 15456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_13
timestamp 1694700623
transform 1 0 2300 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_30
timestamp 1694700623
transform 1 0 3864 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_38
timestamp 1694700623
transform 1 0 4600 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_50
timestamp 1694700623
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_57
timestamp 1694700623
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_65
timestamp 1694700623
transform 1 0 7084 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_73
timestamp 1694700623
transform 1 0 7820 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_94
timestamp 1694700623
transform 1 0 9752 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_106
timestamp 1694700623
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_129
timestamp 1694700623
transform 1 0 12972 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_146
timestamp 1694700623
transform 1 0 14536 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_158
timestamp 1694700623
transform 1 0 15640 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_162
timestamp 1694700623
transform 1 0 16008 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1694700623
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_29
timestamp 1694700623
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_36
timestamp 1694700623
transform 1 0 4416 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_48
timestamp 1694700623
transform 1 0 5520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_79
timestamp 1694700623
transform 1 0 8372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1694700623
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1694700623
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_97
timestamp 1694700623
transform 1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_113
timestamp 1694700623
transform 1 0 11500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_125
timestamp 1694700623
transform 1 0 12604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_137
timestamp 1694700623
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1694700623
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_153
timestamp 1694700623
transform 1 0 15180 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_161
timestamp 1694700623
transform 1 0 15916 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_3
timestamp 1694700623
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_20
timestamp 1694700623
transform 1 0 2944 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_28
timestamp 1694700623
transform 1 0 3680 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_48
timestamp 1694700623
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_70
timestamp 1694700623
transform 1 0 7544 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_78
timestamp 1694700623
transform 1 0 8280 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_91
timestamp 1694700623
transform 1 0 9476 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_95
timestamp 1694700623
transform 1 0 9844 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_102
timestamp 1694700623
transform 1 0 10488 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_106
timestamp 1694700623
transform 1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_118
timestamp 1694700623
transform 1 0 11960 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_126
timestamp 1694700623
transform 1 0 12696 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_136
timestamp 1694700623
transform 1 0 13616 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_148
timestamp 1694700623
transform 1 0 14720 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_160
timestamp 1694700623
transform 1 0 15824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_3
timestamp 1694700623
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_22
timestamp 1694700623
transform 1 0 3128 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_29
timestamp 1694700623
transform 1 0 3772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_33
timestamp 1694700623
transform 1 0 4140 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_41
timestamp 1694700623
transform 1 0 4876 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_49
timestamp 1694700623
transform 1 0 5612 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_58
timestamp 1694700623
transform 1 0 6440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_64
timestamp 1694700623
transform 1 0 6992 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_71
timestamp 1694700623
transform 1 0 7636 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_78
timestamp 1694700623
transform 1 0 8280 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_97
timestamp 1694700623
transform 1 0 10028 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_109
timestamp 1694700623
transform 1 0 11132 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_155
timestamp 1694700623
transform 1 0 15364 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_27
timestamp 1694700623
transform 1 0 3588 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_39
timestamp 1694700623
transform 1 0 4692 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 1694700623
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_74
timestamp 1694700623
transform 1 0 7912 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_79
timestamp 1694700623
transform 1 0 8372 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_89
timestamp 1694700623
transform 1 0 9292 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_101
timestamp 1694700623
transform 1 0 10396 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_109
timestamp 1694700623
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_120
timestamp 1694700623
transform 1 0 12144 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_130
timestamp 1694700623
transform 1 0 13064 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_138
timestamp 1694700623
transform 1 0 13800 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_150
timestamp 1694700623
transform 1 0 14904 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_162
timestamp 1694700623
transform 1 0 16008 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_3
timestamp 1694700623
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_26
timestamp 1694700623
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_29
timestamp 1694700623
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_55
timestamp 1694700623
transform 1 0 6164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_61
timestamp 1694700623
transform 1 0 6716 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_66
timestamp 1694700623
transform 1 0 7176 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_80
timestamp 1694700623
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_85
timestamp 1694700623
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_93
timestamp 1694700623
transform 1 0 9660 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_101
timestamp 1694700623
transform 1 0 10396 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_122
timestamp 1694700623
transform 1 0 12328 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_134
timestamp 1694700623
transform 1 0 13432 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1694700623
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_153
timestamp 1694700623
transform 1 0 15180 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_161
timestamp 1694700623
transform 1 0 15916 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_17
timestamp 1694700623
transform 1 0 2668 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_24
timestamp 1694700623
transform 1 0 3312 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_42
timestamp 1694700623
transform 1 0 4968 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_61
timestamp 1694700623
transform 1 0 6716 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_73
timestamp 1694700623
transform 1 0 7820 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_81
timestamp 1694700623
transform 1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_89
timestamp 1694700623
transform 1 0 9292 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_96
timestamp 1694700623
transform 1 0 9936 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_103
timestamp 1694700623
transform 1 0 10580 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_113
timestamp 1694700623
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_126
timestamp 1694700623
transform 1 0 12696 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_130
timestamp 1694700623
transform 1 0 13064 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_137
timestamp 1694700623
transform 1 0 13708 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_151
timestamp 1694700623
transform 1 0 14996 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_3
timestamp 1694700623
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_16
timestamp 1694700623
transform 1 0 2576 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 1694700623
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_32
timestamp 1694700623
transform 1 0 4048 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_45
timestamp 1694700623
transform 1 0 5244 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_57
timestamp 1694700623
transform 1 0 6348 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_72
timestamp 1694700623
transform 1 0 7728 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1694700623
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_109
timestamp 1694700623
transform 1 0 11132 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_117
timestamp 1694700623
transform 1 0 11868 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_123
timestamp 1694700623
transform 1 0 12420 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_129
timestamp 1694700623
transform 1 0 12972 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_138
timestamp 1694700623
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_141
timestamp 1694700623
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_150
timestamp 1694700623
transform 1 0 14904 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_3
timestamp 1694700623
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_7
timestamp 1694700623
transform 1 0 1748 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_20
timestamp 1694700623
transform 1 0 2944 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_31
timestamp 1694700623
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_43
timestamp 1694700623
transform 1 0 5060 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1694700623
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_69
timestamp 1694700623
transform 1 0 7452 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_81
timestamp 1694700623
transform 1 0 8556 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_87
timestamp 1694700623
transform 1 0 9108 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_106
timestamp 1694700623
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_118
timestamp 1694700623
transform 1 0 11960 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_124
timestamp 1694700623
transform 1 0 12512 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_136
timestamp 1694700623
transform 1 0 13616 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_148
timestamp 1694700623
transform 1 0 14720 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_156
timestamp 1694700623
transform 1 0 15456 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_162
timestamp 1694700623
transform 1 0 16008 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_9
timestamp 1694700623
transform 1 0 1932 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_21
timestamp 1694700623
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1694700623
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_29
timestamp 1694700623
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_37
timestamp 1694700623
transform 1 0 4508 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_50
timestamp 1694700623
transform 1 0 5704 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_66
timestamp 1694700623
transform 1 0 7176 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_71
timestamp 1694700623
transform 1 0 7636 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_81
timestamp 1694700623
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_92
timestamp 1694700623
transform 1 0 9568 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_104
timestamp 1694700623
transform 1 0 10672 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_115
timestamp 1694700623
transform 1 0 11684 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_132
timestamp 1694700623
transform 1 0 13248 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_141
timestamp 1694700623
transform 1 0 14076 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_150
timestamp 1694700623
transform 1 0 14904 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_162
timestamp 1694700623
transform 1 0 16008 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1694700623
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_15
timestamp 1694700623
transform 1 0 2484 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_24
timestamp 1694700623
transform 1 0 3312 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_36
timestamp 1694700623
transform 1 0 4416 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_48
timestamp 1694700623
transform 1 0 5520 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_57
timestamp 1694700623
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_81
timestamp 1694700623
transform 1 0 8556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_85
timestamp 1694700623
transform 1 0 8924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_91
timestamp 1694700623
transform 1 0 9476 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_99
timestamp 1694700623
transform 1 0 10212 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 1694700623
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_118
timestamp 1694700623
transform 1 0 11960 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_126
timestamp 1694700623
transform 1 0 12696 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_161
timestamp 1694700623
transform 1 0 15916 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_9
timestamp 1694700623
transform 1 0 1932 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_21
timestamp 1694700623
transform 1 0 3036 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_26
timestamp 1694700623
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_40
timestamp 1694700623
transform 1 0 4784 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_47
timestamp 1694700623
transform 1 0 5428 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_51
timestamp 1694700623
transform 1 0 5796 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_64
timestamp 1694700623
transform 1 0 6992 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_81
timestamp 1694700623
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_85
timestamp 1694700623
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_102
timestamp 1694700623
transform 1 0 10488 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_114
timestamp 1694700623
transform 1 0 11592 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_127
timestamp 1694700623
transform 1 0 12788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1694700623
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_141
timestamp 1694700623
transform 1 0 14076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_149
timestamp 1694700623
transform 1 0 14812 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_156
timestamp 1694700623
transform 1 0 15456 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_6
timestamp 1694700623
transform 1 0 1656 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_21
timestamp 1694700623
transform 1 0 3036 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_27
timestamp 1694700623
transform 1 0 3588 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_33
timestamp 1694700623
transform 1 0 4140 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_43
timestamp 1694700623
transform 1 0 5060 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_71
timestamp 1694700623
transform 1 0 7636 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_83
timestamp 1694700623
transform 1 0 8740 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_95
timestamp 1694700623
transform 1 0 9844 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_107
timestamp 1694700623
transform 1 0 10948 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1694700623
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_113
timestamp 1694700623
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_121
timestamp 1694700623
transform 1 0 12236 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1694700623
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_149
timestamp 1694700623
transform 1 0 14812 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_6
timestamp 1694700623
transform 1 0 1656 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_18
timestamp 1694700623
transform 1 0 2760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_26
timestamp 1694700623
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1694700623
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1694700623
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_53
timestamp 1694700623
transform 1 0 5980 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_57
timestamp 1694700623
transform 1 0 6348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_77
timestamp 1694700623
transform 1 0 8188 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1694700623
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_88
timestamp 1694700623
transform 1 0 9200 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_100
timestamp 1694700623
transform 1 0 10304 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_111
timestamp 1694700623
transform 1 0 11316 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_125
timestamp 1694700623
transform 1 0 12604 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_138
timestamp 1694700623
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_141
timestamp 1694700623
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_149
timestamp 1694700623
transform 1 0 14812 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_159
timestamp 1694700623
transform 1 0 15732 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1694700623
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_15
timestamp 1694700623
transform 1 0 2484 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_31
timestamp 1694700623
transform 1 0 3956 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_36
timestamp 1694700623
transform 1 0 4416 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_48
timestamp 1694700623
transform 1 0 5520 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1694700623
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_69
timestamp 1694700623
transform 1 0 7452 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_77
timestamp 1694700623
transform 1 0 8188 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_84
timestamp 1694700623
transform 1 0 8832 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_107
timestamp 1694700623
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1694700623
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_116
timestamp 1694700623
transform 1 0 11776 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_128
timestamp 1694700623
transform 1 0 12880 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_140
timestamp 1694700623
transform 1 0 13984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_155
timestamp 1694700623
transform 1 0 15364 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_3
timestamp 1694700623
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_20
timestamp 1694700623
transform 1 0 2944 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_29
timestamp 1694700623
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_42
timestamp 1694700623
transform 1 0 4968 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_58
timestamp 1694700623
transform 1 0 6440 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_70
timestamp 1694700623
transform 1 0 7544 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_79
timestamp 1694700623
transform 1 0 8372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1694700623
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_92
timestamp 1694700623
transform 1 0 9568 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_104
timestamp 1694700623
transform 1 0 10672 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_116
timestamp 1694700623
transform 1 0 11776 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_130
timestamp 1694700623
transform 1 0 13064 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1694700623
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_153
timestamp 1694700623
transform 1 0 15180 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_161
timestamp 1694700623
transform 1 0 15916 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_7
timestamp 1694700623
transform 1 0 1748 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_18
timestamp 1694700623
transform 1 0 2760 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_30
timestamp 1694700623
transform 1 0 3864 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_41
timestamp 1694700623
transform 1 0 4876 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_47
timestamp 1694700623
transform 1 0 5428 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_54
timestamp 1694700623
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_57
timestamp 1694700623
transform 1 0 6348 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_84
timestamp 1694700623
transform 1 0 8832 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_96
timestamp 1694700623
transform 1 0 9936 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_101
timestamp 1694700623
transform 1 0 10396 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_109
timestamp 1694700623
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_120
timestamp 1694700623
transform 1 0 12144 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_139
timestamp 1694700623
transform 1 0 13892 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_143
timestamp 1694700623
transform 1 0 14260 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_151
timestamp 1694700623
transform 1 0 14996 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_6
timestamp 1694700623
transform 1 0 1656 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_15
timestamp 1694700623
transform 1 0 2484 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1694700623
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_47
timestamp 1694700623
transform 1 0 5428 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_55
timestamp 1694700623
transform 1 0 6164 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_62
timestamp 1694700623
transform 1 0 6808 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_72
timestamp 1694700623
transform 1 0 7728 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_76
timestamp 1694700623
transform 1 0 8096 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp 1694700623
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_89
timestamp 1694700623
transform 1 0 9292 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_97
timestamp 1694700623
transform 1 0 10028 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_103
timestamp 1694700623
transform 1 0 10580 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_107
timestamp 1694700623
transform 1 0 10948 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_111
timestamp 1694700623
transform 1 0 11316 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_115
timestamp 1694700623
transform 1 0 11684 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_119
timestamp 1694700623
transform 1 0 12052 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_137
timestamp 1694700623
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_147
timestamp 1694700623
transform 1 0 14628 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_18
timestamp 1694700623
transform 1 0 2760 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_28
timestamp 1694700623
transform 1 0 3680 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_32
timestamp 1694700623
transform 1 0 4048 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_36
timestamp 1694700623
transform 1 0 4416 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_46
timestamp 1694700623
transform 1 0 5336 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_54
timestamp 1694700623
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_57
timestamp 1694700623
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_74
timestamp 1694700623
transform 1 0 7912 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_98
timestamp 1694700623
transform 1 0 10120 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_107
timestamp 1694700623
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1694700623
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1694700623
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1694700623
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 1694700623
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 1694700623
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_161
timestamp 1694700623
transform 1 0 15916 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_7
timestamp 1694700623
transform 1 0 1748 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_22
timestamp 1694700623
transform 1 0 3128 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_55
timestamp 1694700623
transform 1 0 6164 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_63
timestamp 1694700623
transform 1 0 6900 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_71
timestamp 1694700623
transform 1 0 7636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1694700623
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_92
timestamp 1694700623
transform 1 0 9568 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_98
timestamp 1694700623
transform 1 0 10120 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_102
timestamp 1694700623
transform 1 0 10488 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_113
timestamp 1694700623
transform 1 0 11500 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_128
timestamp 1694700623
transform 1 0 12880 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1694700623
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_153
timestamp 1694700623
transform 1 0 15180 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_161
timestamp 1694700623
transform 1 0 15916 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_3
timestamp 1694700623
transform 1 0 1380 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_11
timestamp 1694700623
transform 1 0 2116 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_18
timestamp 1694700623
transform 1 0 2760 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_30
timestamp 1694700623
transform 1 0 3864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_35
timestamp 1694700623
transform 1 0 4324 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_40
timestamp 1694700623
transform 1 0 4784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_52
timestamp 1694700623
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_57
timestamp 1694700623
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_68
timestamp 1694700623
transform 1 0 7360 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_80
timestamp 1694700623
transform 1 0 8464 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_92
timestamp 1694700623
transform 1 0 9568 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_113
timestamp 1694700623
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_121
timestamp 1694700623
transform 1 0 12236 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_145
timestamp 1694700623
transform 1 0 14444 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_157
timestamp 1694700623
transform 1 0 15548 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1694700623
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1694700623
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1694700623
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1694700623
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1694700623
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_53
timestamp 1694700623
transform 1 0 5980 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_64
timestamp 1694700623
transform 1 0 6992 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1694700623
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1694700623
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_85
timestamp 1694700623
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_100
timestamp 1694700623
transform 1 0 10304 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_112
timestamp 1694700623
transform 1 0 11408 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_124
timestamp 1694700623
transform 1 0 12512 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_136
timestamp 1694700623
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1694700623
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_153
timestamp 1694700623
transform 1 0 15180 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1694700623
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1694700623
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1694700623
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_39
timestamp 1694700623
transform 1 0 4692 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_47
timestamp 1694700623
transform 1 0 5428 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_54
timestamp 1694700623
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_64
timestamp 1694700623
transform 1 0 6992 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_72
timestamp 1694700623
transform 1 0 7728 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_84
timestamp 1694700623
transform 1 0 8832 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_96
timestamp 1694700623
transform 1 0 9936 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_101
timestamp 1694700623
transform 1 0 10396 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_109
timestamp 1694700623
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_116
timestamp 1694700623
transform 1 0 11776 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_129
timestamp 1694700623
transform 1 0 12972 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_135
timestamp 1694700623
transform 1 0 13524 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_145
timestamp 1694700623
transform 1 0 14444 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_157
timestamp 1694700623
transform 1 0 15548 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1694700623
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1694700623
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1694700623
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1694700623
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1694700623
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_53
timestamp 1694700623
transform 1 0 5980 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_61
timestamp 1694700623
transform 1 0 6716 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_81
timestamp 1694700623
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_98
timestamp 1694700623
transform 1 0 10120 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_114
timestamp 1694700623
transform 1 0 11592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_134
timestamp 1694700623
transform 1 0 13432 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_148
timestamp 1694700623
transform 1 0 14720 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_160
timestamp 1694700623
transform 1 0 15824 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1694700623
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1694700623
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_27
timestamp 1694700623
transform 1 0 3588 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_29
timestamp 1694700623
transform 1 0 3772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_41
timestamp 1694700623
transform 1 0 4876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_53
timestamp 1694700623
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_57
timestamp 1694700623
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_65
timestamp 1694700623
transform 1 0 7084 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_71
timestamp 1694700623
transform 1 0 7636 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_83
timestamp 1694700623
transform 1 0 8740 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_85
timestamp 1694700623
transform 1 0 8924 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_97
timestamp 1694700623
transform 1 0 10028 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_104
timestamp 1694700623
transform 1 0 10672 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_113
timestamp 1694700623
transform 1 0 11500 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_131
timestamp 1694700623
transform 1 0 13156 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_139
timestamp 1694700623
transform 1 0 13892 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_147
timestamp 1694700623
transform 1 0 14628 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_156
timestamp 1694700623
transform 1 0 15456 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_162
timestamp 1694700623
transform 1 0 16008 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 2576 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1694700623
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  input3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  input4
timestamp 1694700623
transform 1 0 1380 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1694700623
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1694700623
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1694700623
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1694700623
transform 1 0 1932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input10
timestamp 1694700623
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input11
timestamp 1694700623
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input12
timestamp 1694700623
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1694700623
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input14
timestamp 1694700623
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1694700623
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1694700623
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 1694700623
transform -1 0 1932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output18
timestamp 1694700623
transform 1 0 15548 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1694700623
transform 1 0 15732 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output20
timestamp 1694700623
transform 1 0 15548 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 1694700623
transform 1 0 14904 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1694700623
transform 1 0 14076 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  output23
timestamp 1694700623
transform 1 0 12052 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1694700623
transform 1 0 2392 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 1694700623
transform -1 0 1932 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1694700623
transform 1 0 4600 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 1694700623
transform -1 0 8832 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output28
timestamp 1694700623
transform 1 0 12328 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1694700623
transform 1 0 15732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 1694700623
transform 1 0 15548 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1694700623
transform 1 0 15732 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 1694700623
transform 1 0 15548 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_28
timestamp 1694700623
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1694700623
transform -1 0 16376 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_29
timestamp 1694700623
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1694700623
transform -1 0 16376 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_30
timestamp 1694700623
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1694700623
transform -1 0 16376 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_31
timestamp 1694700623
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1694700623
transform -1 0 16376 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_32
timestamp 1694700623
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1694700623
transform -1 0 16376 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_33
timestamp 1694700623
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1694700623
transform -1 0 16376 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_34
timestamp 1694700623
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1694700623
transform -1 0 16376 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_35
timestamp 1694700623
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1694700623
transform -1 0 16376 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_36
timestamp 1694700623
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1694700623
transform -1 0 16376 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_37
timestamp 1694700623
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1694700623
transform -1 0 16376 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_38
timestamp 1694700623
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1694700623
transform -1 0 16376 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_39
timestamp 1694700623
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1694700623
transform -1 0 16376 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_40
timestamp 1694700623
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1694700623
transform -1 0 16376 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_41
timestamp 1694700623
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1694700623
transform -1 0 16376 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_42
timestamp 1694700623
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1694700623
transform -1 0 16376 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_43
timestamp 1694700623
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1694700623
transform -1 0 16376 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_44
timestamp 1694700623
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1694700623
transform -1 0 16376 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_45
timestamp 1694700623
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1694700623
transform -1 0 16376 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_46
timestamp 1694700623
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1694700623
transform -1 0 16376 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_47
timestamp 1694700623
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1694700623
transform -1 0 16376 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_48
timestamp 1694700623
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1694700623
transform -1 0 16376 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_49
timestamp 1694700623
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1694700623
transform -1 0 16376 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_50
timestamp 1694700623
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1694700623
transform -1 0 16376 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_51
timestamp 1694700623
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1694700623
transform -1 0 16376 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_52
timestamp 1694700623
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1694700623
transform -1 0 16376 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_53
timestamp 1694700623
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1694700623
transform -1 0 16376 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_54
timestamp 1694700623
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1694700623
transform -1 0 16376 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_55
timestamp 1694700623
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1694700623
transform -1 0 16376 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 7268 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer2
timestamp 1694700623
transform 1 0 7636 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer3
timestamp 1694700623
transform -1 0 7636 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer4
timestamp 1694700623
transform -1 0 8280 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer5
timestamp 1694700623
transform 1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  rebuffer6
timestamp 1694700623
transform -1 0 8372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer7
timestamp 1694700623
transform -1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer8
timestamp 1694700623
transform 1 0 4140 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer9
timestamp 1694700623
transform 1 0 3680 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  rebuffer10
timestamp 1694700623
transform 1 0 5888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer11
timestamp 1694700623
transform 1 0 6716 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  rebuffer12
timestamp 1694700623
transform -1 0 6716 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  rebuffer13
timestamp 1694700623
transform -1 0 3312 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer14
timestamp 1694700623
transform 1 0 6532 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer15
timestamp 1694700623
transform -1 0 4416 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer16
timestamp 1694700623
transform 1 0 5612 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer17
timestamp 1694700623
transform 1 0 10580 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6348 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6992 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer20
timestamp 1694700623
transform 1 0 6348 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_57
timestamp 1694700623
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_58
timestamp 1694700623
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_59
timestamp 1694700623
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_60
timestamp 1694700623
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_61
timestamp 1694700623
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_62
timestamp 1694700623
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_63
timestamp 1694700623
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_64
timestamp 1694700623
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_65
timestamp 1694700623
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_66
timestamp 1694700623
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_67
timestamp 1694700623
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_68
timestamp 1694700623
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_69
timestamp 1694700623
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_70
timestamp 1694700623
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_71
timestamp 1694700623
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_72
timestamp 1694700623
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_73
timestamp 1694700623
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_74
timestamp 1694700623
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_75
timestamp 1694700623
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_76
timestamp 1694700623
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_77
timestamp 1694700623
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_78
timestamp 1694700623
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_79
timestamp 1694700623
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_80
timestamp 1694700623
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_81
timestamp 1694700623
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_82
timestamp 1694700623
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_83
timestamp 1694700623
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_84
timestamp 1694700623
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_85
timestamp 1694700623
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_86
timestamp 1694700623
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_87
timestamp 1694700623
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_88
timestamp 1694700623
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_89
timestamp 1694700623
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_90
timestamp 1694700623
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_91
timestamp 1694700623
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_92
timestamp 1694700623
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_93
timestamp 1694700623
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_94
timestamp 1694700623
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_95
timestamp 1694700623
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_96
timestamp 1694700623
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_97
timestamp 1694700623
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_98
timestamp 1694700623
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_99
timestamp 1694700623
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_100
timestamp 1694700623
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_101
timestamp 1694700623
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_102
timestamp 1694700623
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_103
timestamp 1694700623
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_104
timestamp 1694700623
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_105
timestamp 1694700623
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_106
timestamp 1694700623
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_107
timestamp 1694700623
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_108
timestamp 1694700623
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_109
timestamp 1694700623
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_110
timestamp 1694700623
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_111
timestamp 1694700623
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_112
timestamp 1694700623
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_113
timestamp 1694700623
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_114
timestamp 1694700623
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_115
timestamp 1694700623
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_116
timestamp 1694700623
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_117
timestamp 1694700623
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_118
timestamp 1694700623
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_119
timestamp 1694700623
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_120
timestamp 1694700623
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_121
timestamp 1694700623
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_122
timestamp 1694700623
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_123
timestamp 1694700623
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_124
timestamp 1694700623
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_125
timestamp 1694700623
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_126
timestamp 1694700623
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_127
timestamp 1694700623
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_128
timestamp 1694700623
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_129
timestamp 1694700623
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_130
timestamp 1694700623
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
<< labels >>
flabel metal4 s 3513 2128 3833 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7331 2128 7651 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 11149 2128 11469 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 14967 2128 15287 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 4580 16424 4900 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 8388 16424 8708 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 12196 16424 12516 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 16004 16424 16324 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2853 2128 3173 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 6671 2128 6991 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 10489 2128 10809 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 14307 2128 14627 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 3920 16424 4240 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 7728 16424 8048 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 11536 16424 11856 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 15344 16424 15664 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 a[0]
port 2 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 a[1]
port 3 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 a[2]
port 4 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 a[3]
port 5 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 a[4]
port 6 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 a[5]
port 7 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 a[6]
port 8 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 a[7]
port 9 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 b[0]
port 10 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 b[1]
port 11 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 b[2]
port 12 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 b[3]
port 13 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 b[4]
port 14 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 b[5]
port 15 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 b[6]
port 16 nsew signal input
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 b[7]
port 17 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 prod[0]
port 18 nsew signal tristate
flabel metal3 s 16699 10888 17499 11008 0 FreeSans 480 0 0 0 prod[10]
port 19 nsew signal tristate
flabel metal3 s 16699 12928 17499 13048 0 FreeSans 480 0 0 0 prod[11]
port 20 nsew signal tristate
flabel metal3 s 16699 14968 17499 15088 0 FreeSans 480 0 0 0 prod[12]
port 21 nsew signal tristate
flabel metal2 s 14830 18843 14886 19643 0 FreeSans 224 90 0 0 prod[13]
port 22 nsew signal tristate
flabel metal2 s 13542 18843 13598 19643 0 FreeSans 224 90 0 0 prod[14]
port 23 nsew signal tristate
flabel metal2 s 12254 18843 12310 19643 0 FreeSans 224 90 0 0 prod[15]
port 24 nsew signal tristate
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 prod[1]
port 25 nsew signal tristate
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 prod[2]
port 26 nsew signal tristate
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 prod[3]
port 27 nsew signal tristate
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 prod[4]
port 28 nsew signal tristate
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 prod[5]
port 29 nsew signal tristate
flabel metal3 s 16699 3408 17499 3528 0 FreeSans 480 0 0 0 prod[6]
port 30 nsew signal tristate
flabel metal3 s 16699 5448 17499 5568 0 FreeSans 480 0 0 0 prod[7]
port 31 nsew signal tristate
flabel metal3 s 16699 7488 17499 7608 0 FreeSans 480 0 0 0 prod[8]
port 32 nsew signal tristate
flabel metal3 s 16699 9528 17499 9648 0 FreeSans 480 0 0 0 prod[9]
port 33 nsew signal tristate
rlabel metal1 8740 17408 8740 17408 0 VGND
rlabel metal1 8740 16864 8740 16864 0 VPWR
rlabel metal1 6532 4794 6532 4794 0 _000_
rlabel metal1 7452 4522 7452 4522 0 _001_
rlabel metal1 7682 4590 7682 4590 0 _002_
rlabel metal1 7912 4658 7912 4658 0 _003_
rlabel metal1 8234 4046 8234 4046 0 _004_
rlabel metal1 9292 3706 9292 3706 0 _005_
rlabel metal1 10488 2414 10488 2414 0 _006_
rlabel metal1 11178 2958 11178 2958 0 _007_
rlabel metal1 10718 2618 10718 2618 0 _008_
rlabel metal1 14306 3468 14306 3468 0 _009_
rlabel metal1 1886 12614 1886 12614 0 _010_
rlabel metal1 6026 10676 6026 10676 0 _011_
rlabel metal1 5198 9010 5198 9010 0 _012_
rlabel metal1 4324 9622 4324 9622 0 _013_
rlabel metal1 3450 9554 3450 9554 0 _014_
rlabel metal1 3864 9554 3864 9554 0 _015_
rlabel metal1 13294 3502 13294 3502 0 _016_
rlabel metal1 9660 3570 9660 3570 0 _017_
rlabel metal1 12558 4046 12558 4046 0 _018_
rlabel metal2 8970 7922 8970 7922 0 _019_
rlabel metal1 9338 5780 9338 5780 0 _020_
rlabel metal1 10212 5678 10212 5678 0 _021_
rlabel metal1 8418 6766 8418 6766 0 _022_
rlabel metal1 8497 6426 8497 6426 0 _023_
rlabel metal1 12006 6290 12006 6290 0 _024_
rlabel metal2 11546 5542 11546 5542 0 _025_
rlabel metal1 11960 4114 11960 4114 0 _026_
rlabel metal1 11270 4590 11270 4590 0 _027_
rlabel metal2 10074 5678 10074 5678 0 _028_
rlabel metal1 9844 5202 9844 5202 0 _029_
rlabel metal1 10442 4726 10442 4726 0 _030_
rlabel metal1 11316 4114 11316 4114 0 _031_
rlabel metal2 12650 3740 12650 3740 0 _032_
rlabel metal1 13708 3570 13708 3570 0 _033_
rlabel metal1 13984 3706 13984 3706 0 _034_
rlabel metal1 14306 4080 14306 4080 0 _035_
rlabel metal1 14858 5678 14858 5678 0 _036_
rlabel metal1 2346 14790 2346 14790 0 _037_
rlabel metal1 2024 13974 2024 13974 0 _038_
rlabel metal1 1932 13362 1932 13362 0 _039_
rlabel metal1 2484 10710 2484 10710 0 _040_
rlabel metal1 4922 10098 4922 10098 0 _041_
rlabel metal1 6716 11050 6716 11050 0 _042_
rlabel metal1 6256 10234 6256 10234 0 _043_
rlabel metal1 5520 10642 5520 10642 0 _044_
rlabel metal1 5658 12274 5658 12274 0 _045_
rlabel metal1 5198 10064 5198 10064 0 _046_
rlabel metal1 2162 10540 2162 10540 0 _047_
rlabel metal2 2438 10404 2438 10404 0 _048_
rlabel metal1 3910 10472 3910 10472 0 _049_
rlabel metal1 4232 10030 4232 10030 0 _050_
rlabel metal1 14122 5678 14122 5678 0 _051_
rlabel metal1 12696 4114 12696 4114 0 _052_
rlabel metal1 13018 5678 13018 5678 0 _053_
rlabel metal1 11776 5678 11776 5678 0 _054_
rlabel metal1 11546 5644 11546 5644 0 _055_
rlabel metal1 8234 7310 8234 7310 0 _056_
rlabel metal1 8602 7446 8602 7446 0 _057_
rlabel metal1 10810 7446 10810 7446 0 _058_
rlabel metal1 9246 7446 9246 7446 0 _059_
rlabel metal1 9246 7820 9246 7820 0 _060_
rlabel metal1 8004 9350 8004 9350 0 _061_
rlabel metal2 9706 8160 9706 8160 0 _062_
rlabel metal1 9062 6698 9062 6698 0 _063_
rlabel metal1 10350 7480 10350 7480 0 _064_
rlabel metal2 10166 7174 10166 7174 0 _065_
rlabel metal1 10488 7174 10488 7174 0 _066_
rlabel metal1 11684 6630 11684 6630 0 _067_
rlabel metal1 12374 5814 12374 5814 0 _068_
rlabel metal2 13202 5372 13202 5372 0 _069_
rlabel metal1 12834 5882 12834 5882 0 _070_
rlabel metal1 13340 5338 13340 5338 0 _071_
rlabel metal1 14030 5746 14030 5746 0 _072_
rlabel metal2 14674 6086 14674 6086 0 _073_
rlabel metal1 14674 6256 14674 6256 0 _074_
rlabel metal1 14812 6426 14812 6426 0 _075_
rlabel metal1 4232 10574 4232 10574 0 _076_
rlabel metal2 2714 13396 2714 13396 0 _077_
rlabel metal1 2346 12274 2346 12274 0 _078_
rlabel metal1 3174 12206 3174 12206 0 _079_
rlabel metal1 6026 13294 6026 13294 0 _080_
rlabel metal1 6026 12274 6026 12274 0 _081_
rlabel metal1 4278 12138 4278 12138 0 _082_
rlabel metal1 3450 11662 3450 11662 0 _083_
rlabel metal1 3864 12070 3864 12070 0 _084_
rlabel metal1 3818 10642 3818 10642 0 _085_
rlabel metal2 4186 11968 4186 11968 0 _086_
rlabel metal1 4554 10064 4554 10064 0 _087_
rlabel metal1 10810 11016 10810 11016 0 _088_
rlabel metal1 10856 11118 10856 11118 0 _089_
rlabel metal1 11224 11186 11224 11186 0 _090_
rlabel viali 11914 11110 11914 11110 0 _091_
rlabel metal1 14168 7854 14168 7854 0 _092_
rlabel metal1 13156 7242 13156 7242 0 _093_
rlabel metal1 11822 7446 11822 7446 0 _094_
rlabel metal1 12006 6766 12006 6766 0 _095_
rlabel metal1 12144 6970 12144 6970 0 _096_
rlabel metal1 7590 9554 7590 9554 0 _097_
rlabel metal1 7774 9486 7774 9486 0 _098_
rlabel metal1 8372 8942 8372 8942 0 _099_
rlabel metal1 11454 8976 11454 8976 0 _100_
rlabel metal1 8372 12886 8372 12886 0 _101_
rlabel metal1 10166 8398 10166 8398 0 _102_
rlabel metal1 11730 8398 11730 8398 0 _103_
rlabel metal1 12466 8908 12466 8908 0 _104_
rlabel metal1 12006 8466 12006 8466 0 _105_
rlabel metal2 12466 8058 12466 8058 0 _106_
rlabel metal1 12742 7922 12742 7922 0 _107_
rlabel metal1 12788 7514 12788 7514 0 _108_
rlabel metal1 13064 7922 13064 7922 0 _109_
rlabel metal1 14076 7922 14076 7922 0 _110_
rlabel metal1 14858 8058 14858 8058 0 _111_
rlabel metal1 14904 7514 14904 7514 0 _112_
rlabel metal1 15456 9554 15456 9554 0 _113_
rlabel metal1 9752 11730 9752 11730 0 _114_
rlabel metal1 8740 11186 8740 11186 0 _115_
rlabel metal1 9154 11730 9154 11730 0 _116_
rlabel metal1 10074 11764 10074 11764 0 _117_
rlabel metal1 5612 13294 5612 13294 0 _118_
rlabel metal1 4186 14314 4186 14314 0 _119_
rlabel metal1 3174 13702 3174 13702 0 _120_
rlabel metal1 3542 14382 3542 14382 0 _121_
rlabel metal1 3358 14416 3358 14416 0 _122_
rlabel via1 4278 14450 4278 14450 0 _123_
rlabel metal1 3818 13906 3818 13906 0 _124_
rlabel metal1 4646 13294 4646 13294 0 _125_
rlabel metal1 4646 12852 4646 12852 0 _126_
rlabel metal1 5336 13906 5336 13906 0 _127_
rlabel metal1 4508 12614 4508 12614 0 _128_
rlabel metal1 5152 13906 5152 13906 0 _129_
rlabel metal1 4462 11866 4462 11866 0 _130_
rlabel metal1 10074 11662 10074 11662 0 _131_
rlabel metal1 10994 11730 10994 11730 0 _132_
rlabel metal1 11822 11866 11822 11866 0 _133_
rlabel metal1 12190 11220 12190 11220 0 _134_
rlabel metal1 14444 9554 14444 9554 0 _135_
rlabel metal1 13708 9554 13708 9554 0 _136_
rlabel via1 10534 9469 10534 9469 0 _137_
rlabel metal1 8004 9622 8004 9622 0 _138_
rlabel metal1 8924 10234 8924 10234 0 _139_
rlabel metal1 8480 9962 8480 9962 0 _140_
rlabel metal1 9430 9962 9430 9962 0 _141_
rlabel metal1 10442 9520 10442 9520 0 _142_
rlabel metal1 12558 9996 12558 9996 0 _143_
rlabel metal1 11454 9554 11454 9554 0 _144_
rlabel metal1 12098 9010 12098 9010 0 _145_
rlabel metal1 12650 9928 12650 9928 0 _146_
rlabel metal1 13018 8908 13018 8908 0 _147_
rlabel metal1 13386 9554 13386 9554 0 _148_
rlabel metal1 14674 9486 14674 9486 0 _149_
rlabel metal1 15410 9486 15410 9486 0 _150_
rlabel metal2 14858 9588 14858 9588 0 _151_
rlabel metal1 15088 11118 15088 11118 0 _152_
rlabel metal1 11408 12206 11408 12206 0 _153_
rlabel metal1 8894 12886 8894 12886 0 _154_
rlabel metal1 8924 11866 8924 11866 0 _155_
rlabel metal1 10350 12784 10350 12784 0 _156_
rlabel metal1 7398 13158 7398 13158 0 _157_
rlabel metal1 10902 13260 10902 13260 0 _158_
rlabel metal1 10534 12954 10534 12954 0 _159_
rlabel metal1 11454 13328 11454 13328 0 _160_
rlabel metal2 3818 14688 3818 14688 0 _161_
rlabel metal1 4738 15028 4738 15028 0 _162_
rlabel metal2 5198 14586 5198 14586 0 _163_
rlabel metal1 5528 14246 5528 14246 0 _164_
rlabel metal1 5612 14042 5612 14042 0 _165_
rlabel metal1 11638 13362 11638 13362 0 _166_
rlabel metal1 12144 12206 12144 12206 0 _167_
rlabel metal1 13018 12308 13018 12308 0 _168_
rlabel metal1 12834 12138 12834 12138 0 _169_
rlabel metal1 13662 11730 13662 11730 0 _170_
rlabel metal1 13478 10608 13478 10608 0 _171_
rlabel metal1 10074 10030 10074 10030 0 _172_
rlabel metal1 9752 10098 9752 10098 0 _173_
rlabel metal1 12190 10064 12190 10064 0 _174_
rlabel metal1 12788 10710 12788 10710 0 _175_
rlabel metal2 12742 10438 12742 10438 0 _176_
rlabel metal1 13662 10676 13662 10676 0 _177_
rlabel metal1 14582 11152 14582 11152 0 _178_
rlabel metal1 15318 11696 15318 11696 0 _179_
rlabel metal1 14904 11322 14904 11322 0 _180_
rlabel metal1 14720 12818 14720 12818 0 _181_
rlabel metal1 12742 13362 12742 13362 0 _182_
rlabel metal1 7728 14314 7728 14314 0 _183_
rlabel metal1 6992 14314 6992 14314 0 _184_
rlabel metal1 9890 14280 9890 14280 0 _185_
rlabel metal1 8648 13226 8648 13226 0 _186_
rlabel metal1 8372 13838 8372 13838 0 _187_
rlabel metal1 8288 13158 8288 13158 0 _188_
rlabel metal1 8648 13838 8648 13838 0 _189_
rlabel metal1 9108 13906 9108 13906 0 _190_
rlabel metal1 9568 14042 9568 14042 0 _191_
rlabel metal1 10396 13906 10396 13906 0 _192_
rlabel metal1 10672 14790 10672 14790 0 _193_
rlabel metal2 10902 14178 10902 14178 0 _194_
rlabel metal1 11684 14382 11684 14382 0 _195_
rlabel metal1 12466 14552 12466 14552 0 _196_
rlabel metal2 12742 13770 12742 13770 0 _197_
rlabel metal1 13156 14790 13156 14790 0 _198_
rlabel metal1 13478 13260 13478 13260 0 _199_
rlabel metal1 13708 12342 13708 12342 0 _200_
rlabel metal1 13202 10472 13202 10472 0 _201_
rlabel metal1 9936 10166 9936 10166 0 _202_
rlabel metal2 13478 11458 13478 11458 0 _203_
rlabel metal1 14168 12750 14168 12750 0 _204_
rlabel metal1 14122 13294 14122 13294 0 _205_
rlabel metal1 13846 14994 13846 14994 0 _206_
rlabel metal1 12834 14892 12834 14892 0 _207_
rlabel metal1 10212 14994 10212 14994 0 _208_
rlabel metal1 7452 15674 7452 15674 0 _209_
rlabel metal1 6992 14926 6992 14926 0 _210_
rlabel metal1 8648 15538 8648 15538 0 _211_
rlabel metal1 8832 13838 8832 13838 0 _212_
rlabel metal1 9384 15470 9384 15470 0 _213_
rlabel metal1 10212 16082 10212 16082 0 _214_
rlabel metal1 9706 15402 9706 15402 0 _215_
rlabel metal1 10212 15062 10212 15062 0 _216_
rlabel metal1 10350 14790 10350 14790 0 _217_
rlabel metal1 10994 15096 10994 15096 0 _218_
rlabel metal1 12466 15062 12466 15062 0 _219_
rlabel metal1 12880 16218 12880 16218 0 _220_
rlabel metal1 14352 14994 14352 14994 0 _221_
rlabel metal1 13938 14926 13938 14926 0 _222_
rlabel metal1 9062 16558 9062 16558 0 _223_
rlabel metal1 6440 15946 6440 15946 0 _224_
rlabel metal1 6670 16558 6670 16558 0 _225_
rlabel metal1 6670 15130 6670 15130 0 _226_
rlabel metal1 2484 7854 2484 7854 0 _227_
rlabel metal1 7268 16558 7268 16558 0 _228_
rlabel metal2 7222 16966 7222 16966 0 _229_
rlabel metal1 9062 16694 9062 16694 0 _230_
rlabel metal1 10258 16592 10258 16592 0 _231_
rlabel metal2 10350 16915 10350 16915 0 _232_
rlabel metal1 11086 16558 11086 16558 0 _233_
rlabel metal1 12926 16048 12926 16048 0 _234_
rlabel metal2 14398 16286 14398 16286 0 _235_
rlabel metal1 13340 16558 13340 16558 0 _236_
rlabel metal1 10258 16694 10258 16694 0 _237_
rlabel metal1 7406 16524 7406 16524 0 _238_
rlabel metal1 7774 16626 7774 16626 0 _239_
rlabel metal1 10626 17136 10626 17136 0 _240_
rlabel metal1 11684 16082 11684 16082 0 _241_
rlabel metal1 11316 16082 11316 16082 0 _242_
rlabel metal1 12535 16150 12535 16150 0 _243_
rlabel metal1 13110 17136 13110 17136 0 _244_
rlabel metal1 12742 15946 12742 15946 0 _245_
rlabel metal2 12926 16796 12926 16796 0 _246_
rlabel metal1 2484 7378 2484 7378 0 _247_
rlabel metal2 12650 16796 12650 16796 0 _248_
rlabel metal1 12650 16218 12650 16218 0 _249_
rlabel metal2 8602 3094 8602 3094 0 _250_
rlabel metal2 2438 7888 2438 7888 0 _251_
rlabel metal1 3542 2958 3542 2958 0 _252_
rlabel metal1 2162 12750 2162 12750 0 _253_
rlabel metal1 2070 13260 2070 13260 0 _254_
rlabel metal1 1978 7854 1978 7854 0 _255_
rlabel metal1 2254 7514 2254 7514 0 _256_
rlabel viali 3918 7377 3918 7377 0 _257_
rlabel metal1 4048 8262 4048 8262 0 _258_
rlabel metal1 3266 7718 3266 7718 0 _259_
rlabel metal1 2576 8058 2576 8058 0 _260_
rlabel metal1 7406 9690 7406 9690 0 _261_
rlabel metal1 4554 7174 4554 7174 0 _262_
rlabel metal1 4600 7378 4600 7378 0 _263_
rlabel metal1 3588 7854 3588 7854 0 _264_
rlabel metal1 7360 3026 7360 3026 0 _265_
rlabel metal1 7544 7446 7544 7446 0 _266_
rlabel metal1 4324 5610 4324 5610 0 _267_
rlabel metal1 4922 6766 4922 6766 0 _268_
rlabel metal1 3680 4182 3680 4182 0 _269_
rlabel metal1 9154 10030 9154 10030 0 _270_
rlabel metal1 3772 4114 3772 4114 0 _271_
rlabel metal1 2576 14382 2576 14382 0 _272_
rlabel metal2 2622 5440 2622 5440 0 _273_
rlabel metal1 2208 4590 2208 4590 0 _274_
rlabel metal1 2484 4590 2484 4590 0 _275_
rlabel metal2 2806 4420 2806 4420 0 _276_
rlabel metal1 2668 4114 2668 4114 0 _277_
rlabel metal1 3174 3026 3174 3026 0 _278_
rlabel metal1 4462 2992 4462 2992 0 _279_
rlabel metal1 5842 2924 5842 2924 0 _280_
rlabel via1 4555 5678 4555 5678 0 _281_
rlabel metal2 5106 5916 5106 5916 0 _282_
rlabel metal1 5290 3026 5290 3026 0 _283_
rlabel metal1 4186 4556 4186 4556 0 _284_
rlabel metal1 4324 5202 4324 5202 0 _285_
rlabel metal1 5842 3536 5842 3536 0 _286_
rlabel metal1 5658 2890 5658 2890 0 _287_
rlabel metal1 7222 3128 7222 3128 0 _288_
rlabel metal2 8510 2652 8510 2652 0 _289_
rlabel metal1 7774 2448 7774 2448 0 _290_
rlabel metal1 7682 3026 7682 3026 0 _291_
rlabel metal1 8786 3094 8786 3094 0 _292_
rlabel metal1 11454 3026 11454 3026 0 _293_
rlabel metal1 6348 8534 6348 8534 0 _294_
rlabel metal1 6302 8602 6302 8602 0 _295_
rlabel metal1 7130 8840 7130 8840 0 _296_
rlabel metal1 10166 2414 10166 2414 0 _297_
rlabel metal1 9200 3026 9200 3026 0 _298_
rlabel metal1 8464 5202 8464 5202 0 _299_
rlabel metal1 9200 5066 9200 5066 0 _300_
rlabel metal1 8694 8058 8694 8058 0 _301_
rlabel metal1 8878 5100 8878 5100 0 _302_
rlabel metal1 8878 4114 8878 4114 0 _303_
rlabel metal1 5934 3468 5934 3468 0 _304_
rlabel metal1 6164 3502 6164 3502 0 _305_
rlabel metal1 7222 4114 7222 4114 0 _306_
rlabel metal1 4922 4658 4922 4658 0 _307_
rlabel metal1 5152 6290 5152 6290 0 _308_
rlabel metal1 6302 7514 6302 7514 0 _309_
rlabel metal1 6302 6426 6302 6426 0 _310_
rlabel metal1 5658 6630 5658 6630 0 _311_
rlabel metal1 5950 6358 5950 6358 0 _312_
rlabel metal1 5888 5746 5888 5746 0 _313_
rlabel metal2 2806 5729 2806 5729 0 a[0]
rlabel metal3 820 7548 820 7548 0 a[1]
rlabel metal3 820 2788 820 2788 0 a[2]
rlabel metal3 820 5508 820 5508 0 a[3]
rlabel metal2 7774 1520 7774 1520 0 a[4]
rlabel metal2 9062 1027 9062 1027 0 a[5]
rlabel metal2 7130 1027 7130 1027 0 a[6]
rlabel metal3 820 10268 820 10268 0 a[7]
rlabel metal3 866 4148 866 4148 0 b[0]
rlabel metal3 843 4828 843 4828 0 b[1]
rlabel metal3 820 3468 820 3468 0 b[2]
rlabel metal3 820 6868 820 6868 0 b[3]
rlabel metal3 1050 10948 1050 10948 0 b[4]
rlabel metal3 1050 12308 1050 12308 0 b[5]
rlabel metal3 820 12988 820 12988 0 b[6]
rlabel metal3 820 14348 820 14348 0 b[7]
rlabel metal1 3266 5678 3266 5678 0 net1
rlabel metal1 1794 5202 1794 5202 0 net10
rlabel metal1 3588 6290 3588 6290 0 net11
rlabel metal2 1702 6052 1702 6052 0 net12
rlabel metal1 5888 10030 5888 10030 0 net13
rlabel metal1 6302 9010 6302 9010 0 net14
rlabel metal1 2346 13192 2346 13192 0 net15
rlabel metal2 2300 13906 2300 13906 0 net16
rlabel metal1 1748 8058 1748 8058 0 net17
rlabel metal2 15686 10948 15686 10948 0 net18
rlabel metal1 15364 12750 15364 12750 0 net19
rlabel metal1 4784 7378 4784 7378 0 net2
rlabel metal2 14122 15164 14122 15164 0 net20
rlabel metal1 14812 16762 14812 16762 0 net21
rlabel metal1 13800 16762 13800 16762 0 net22
rlabel metal2 12190 16966 12190 16966 0 net23
rlabel metal1 2438 8466 2438 8466 0 net24
rlabel metal1 2277 10030 2277 10030 0 net25
rlabel metal1 4554 2414 4554 2414 0 net26
rlabel metal1 8648 2414 8648 2414 0 net27
rlabel metal2 12466 2652 12466 2652 0 net28
rlabel metal1 15226 3502 15226 3502 0 net29
rlabel metal2 1978 4318 1978 4318 0 net3
rlabel metal1 15686 5712 15686 5712 0 net30
rlabel metal1 15778 7888 15778 7888 0 net31
rlabel metal1 15778 9486 15778 9486 0 net32
rlabel metal1 6118 4658 6118 4658 0 net33
rlabel metal1 7544 5678 7544 5678 0 net34
rlabel metal1 8004 5678 8004 5678 0 net35
rlabel metal1 8188 3502 8188 3502 0 net36
rlabel metal2 7038 3264 7038 3264 0 net37
rlabel metal1 7682 5168 7682 5168 0 net38
rlabel metal1 4462 7412 4462 7412 0 net39
rlabel metal2 1794 5134 1794 5134 0 net4
rlabel metal1 3726 3060 3726 3060 0 net40
rlabel metal1 2070 7480 2070 7480 0 net41
rlabel metal2 6118 8500 6118 8500 0 net42
rlabel metal1 6578 9962 6578 9962 0 net43
rlabel metal1 6624 13294 6624 13294 0 net44
rlabel metal2 2806 13634 2806 13634 0 net45
rlabel metal1 6256 12954 6256 12954 0 net46
rlabel metal1 4278 4114 4278 4114 0 net47
rlabel metal1 5474 2958 5474 2958 0 net48
rlabel metal1 10534 4658 10534 4658 0 net49
rlabel metal1 8004 6766 8004 6766 0 net5
rlabel metal1 7084 5202 7084 5202 0 net50
rlabel metal1 6762 10574 6762 10574 0 net51
rlabel metal1 6072 12206 6072 12206 0 net52
rlabel viali 9423 5204 9423 5204 0 net6
rlabel metal1 7268 2618 7268 2618 0 net7
rlabel metal2 7314 8092 7314 8092 0 net8
rlabel metal1 1610 5610 1610 5610 0 net9
rlabel metal3 820 8908 820 8908 0 prod[0]
rlabel metal1 16008 10778 16008 10778 0 prod[10]
rlabel metal2 15962 13073 15962 13073 0 prod[11]
rlabel metal1 16008 15334 16008 15334 0 prod[12]
rlabel metal1 15088 17306 15088 17306 0 prod[13]
rlabel metal1 14076 17306 14076 17306 0 prod[14]
rlabel metal1 12512 17238 12512 17238 0 prod[15]
rlabel metal3 1694 8228 1694 8228 0 prod[1]
rlabel metal3 1096 9588 1096 9588 0 prod[2]
rlabel metal2 4554 1520 4554 1520 0 prod[3]
rlabel metal2 8418 1520 8418 1520 0 prod[4]
rlabel metal2 12282 1571 12282 1571 0 prod[5]
rlabel metal2 15962 3553 15962 3553 0 prod[6]
rlabel metal1 16008 5542 16008 5542 0 prod[7]
rlabel metal2 15962 7633 15962 7633 0 prod[8]
rlabel metal1 16008 9894 16008 9894 0 prod[9]
<< properties >>
string FIXED_BBOX 0 0 17499 19643
<< end >>
