magic
tech sky130A
magscale 1 2
timestamp 1699032937
<< obsli1 >>
rect 1104 2159 16376 17425
<< obsm1 >>
rect 934 2128 16376 17456
<< metal2 >>
rect 12254 18843 12310 19643
rect 13542 18843 13598 19643
rect 14830 18843 14886 19643
rect 4526 0 4582 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 12254 0 12310 800
<< obsm2 >>
rect 938 18787 12198 18986
rect 12366 18787 13486 18986
rect 13654 18787 14774 18986
rect 14942 18787 16082 18986
rect 938 856 16082 18787
rect 938 800 4470 856
rect 4638 800 7046 856
rect 7214 800 7690 856
rect 7858 800 8334 856
rect 8502 800 8978 856
rect 9146 800 12198 856
rect 12366 800 16082 856
<< metal3 >>
rect 16699 14968 17499 15088
rect 0 14288 800 14408
rect 0 12928 800 13048
rect 16699 12928 17499 13048
rect 0 12248 800 12368
rect 0 10888 800 11008
rect 16699 10888 17499 11008
rect 0 10208 800 10328
rect 0 9528 800 9648
rect 16699 9528 17499 9648
rect 0 8848 800 8968
rect 0 8168 800 8288
rect 0 7488 800 7608
rect 16699 7488 17499 7608
rect 0 6808 800 6928
rect 0 6128 800 6248
rect 0 5448 800 5568
rect 16699 5448 17499 5568
rect 0 4768 800 4888
rect 0 4088 800 4208
rect 0 3408 800 3528
rect 16699 3408 17499 3528
rect 0 2728 800 2848
<< obsm3 >>
rect 800 15168 16699 17441
rect 800 14888 16619 15168
rect 800 14488 16699 14888
rect 880 14208 16699 14488
rect 800 13128 16699 14208
rect 880 12848 16619 13128
rect 800 12448 16699 12848
rect 880 12168 16699 12448
rect 800 11088 16699 12168
rect 880 10808 16619 11088
rect 800 10408 16699 10808
rect 880 10128 16699 10408
rect 800 9728 16699 10128
rect 880 9448 16619 9728
rect 800 9048 16699 9448
rect 880 8768 16699 9048
rect 800 8368 16699 8768
rect 880 8088 16699 8368
rect 800 7688 16699 8088
rect 880 7408 16619 7688
rect 800 7008 16699 7408
rect 880 6728 16699 7008
rect 800 6328 16699 6728
rect 880 6048 16699 6328
rect 800 5648 16699 6048
rect 880 5368 16619 5648
rect 800 4968 16699 5368
rect 880 4688 16699 4968
rect 800 4288 16699 4688
rect 880 4008 16699 4288
rect 800 3608 16699 4008
rect 880 3328 16619 3608
rect 800 2928 16699 3328
rect 880 2648 16699 2928
rect 800 2143 16699 2648
<< metal4 >>
rect 2853 2128 3173 17456
rect 3513 2128 3833 17456
rect 6671 2128 6991 17456
rect 7331 2128 7651 17456
rect 10489 2128 10809 17456
rect 11149 2128 11469 17456
rect 14307 2128 14627 17456
rect 14967 2128 15287 17456
<< metal5 >>
rect 1056 16004 16424 16324
rect 1056 15344 16424 15664
rect 1056 12196 16424 12516
rect 1056 11536 16424 11856
rect 1056 8388 16424 8708
rect 1056 7728 16424 8048
rect 1056 4580 16424 4900
rect 1056 3920 16424 4240
<< labels >>
rlabel metal4 s 3513 2128 3833 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 7331 2128 7651 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 11149 2128 11469 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 14967 2128 15287 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 4580 16424 4900 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 8388 16424 8708 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 12196 16424 12516 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 16004 16424 16324 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 2853 2128 3173 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 6671 2128 6991 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 10489 2128 10809 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 14307 2128 14627 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 3920 16424 4240 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 7728 16424 8048 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 11536 16424 11856 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 15344 16424 15664 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 6128 800 6248 6 a[0]
port 3 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 a[1]
port 4 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 a[2]
port 5 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 a[3]
port 6 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 a[4]
port 7 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 a[5]
port 8 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 a[6]
port 9 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 a[7]
port 10 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 b[0]
port 11 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 b[1]
port 12 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 b[2]
port 13 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 b[3]
port 14 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 b[4]
port 15 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 b[5]
port 16 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 b[6]
port 17 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 b[7]
port 18 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 prod[0]
port 19 nsew signal output
rlabel metal3 s 16699 10888 17499 11008 6 prod[10]
port 20 nsew signal output
rlabel metal3 s 16699 12928 17499 13048 6 prod[11]
port 21 nsew signal output
rlabel metal3 s 16699 14968 17499 15088 6 prod[12]
port 22 nsew signal output
rlabel metal2 s 14830 18843 14886 19643 6 prod[13]
port 23 nsew signal output
rlabel metal2 s 13542 18843 13598 19643 6 prod[14]
port 24 nsew signal output
rlabel metal2 s 12254 18843 12310 19643 6 prod[15]
port 25 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 prod[1]
port 26 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 prod[2]
port 27 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 prod[3]
port 28 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 prod[4]
port 29 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 prod[5]
port 30 nsew signal output
rlabel metal3 s 16699 3408 17499 3528 6 prod[6]
port 31 nsew signal output
rlabel metal3 s 16699 5448 17499 5568 6 prod[7]
port 32 nsew signal output
rlabel metal3 s 16699 7488 17499 7608 6 prod[8]
port 33 nsew signal output
rlabel metal3 s 16699 9528 17499 9648 6 prod[9]
port 34 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 17499 19643
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1215972
string GDS_FILE /openlane/openlane/pes_vedic_mul/runs/run_4/results/signoff/pes_vedic_mul.magic.gds
string GDS_START 331526
<< end >>

