* NGSPICE file created from pes_vedic_mul.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

.subckt pes_vedic_mul VGND VPWR a[0] a[1] a[2] a[3] a[4] a[5] a[6] a[7] b[0] b[1]
+ b[2] b[3] b[4] b[5] b[6] b[7] prod[0] prod[10] prod[11] prod[12] prod[13] prod[14]
+ prod[15] prod[1] prod[2] prod[3] prod[4] prod[5] prod[6] prod[7] prod[8] prod[9]
XFILLER_0_27_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_432_ _121_ _162_ _164_ VGND VGND VPWR VPWR _196_ sky130_fd_sc_hd__and3_1
X_363_ _126_ _127_ VGND VGND VPWR VPWR _128_ sky130_fd_sc_hd__nand2_1
X_501_ _247_ net2 VGND VGND VPWR VPWR _251_ sky130_fd_sc_hd__nand2_1
Xrebuffer7 _264_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_415_ _152_ _179_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__xor2_1
X_346_ _092_ _110_ VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_329_ _058_ _066_ VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_8_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_594_ _272_ _270_ _281_ _313_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__a31o_1
Xrebuffer17 _027_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_27_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput20 net20 VGND VGND VPWR VPWR prod[12] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_18_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_577_ _254_ net14 _294_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput31 net31 VGND VGND VPWR VPWR prod[8] sky130_fd_sc_hd__buf_2
XFILLER_0_27_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_431_ _193_ _194_ VGND VGND VPWR VPWR _195_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_21_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_362_ _080_ _125_ _118_ VGND VGND VPWR VPWR _127_ sky130_fd_sc_hd__nand3_1
Xrebuffer8 _264_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
X_500_ net10 VGND VGND VPWR VPWR _247_ sky130_fd_sc_hd__buf_6
XFILLER_0_13_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_629_ _059_ _062_ _063_ VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_20_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_414_ _170_ _178_ VGND VGND VPWR VPWR _179_ sky130_fd_sc_hd__xor2_1
X_345_ _093_ _109_ VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_328_ _053_ _070_ _069_ VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_9_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_24_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_84 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer18 _313_ VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_593_ _272_ _270_ _313_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_27_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput21 net21 VGND VGND VPWR VPWR prod[13] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_18_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput32 net32 VGND VGND VPWR VPWR prod[9] sky130_fd_sc_hd__clkbuf_4
X_576_ net42 net13 VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__nand2_2
XFILLER_0_5_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_430_ _158_ _192_ VGND VGND VPWR VPWR _194_ sky130_fd_sc_hd__nand2_1
X_361_ _080_ _118_ _125_ VGND VGND VPWR VPWR _126_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_9 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer9 _257_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_1
X_628_ _019_ _299_ _300_ VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__a21oi_1
X_559_ net4 VGND VGND VPWR VPWR _308_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_413_ _171_ _177_ VGND VGND VPWR VPWR _178_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_8_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_344_ _107_ _108_ VGND VGND VPWR VPWR _109_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_327_ _090_ _091_ VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_592_ _306_ _003_ _001_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer19 _308_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dlygate4sd1_1
Xoutput22 net22 VGND VGND VPWR VPWR prod[14] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_27_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_575_ _253_ net15 VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_360_ _123_ _124_ VGND VGND VPWR VPWR _125_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_489_ _292_ _007_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__xnor2_1
X_558_ _284_ _285_ _273_ VGND VGND VPWR VPWR _307_ sky130_fd_sc_hd__a21boi_1
X_627_ _060_ _061_ _019_ VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__or3_4
X_412_ _175_ _176_ VGND VGND VPWR VPWR _177_ sky130_fd_sc_hd__and2_1
X_343_ _094_ _096_ _106_ VGND VGND VPWR VPWR _108_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_326_ _088_ _089_ VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_591_ _024_ _025_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__or2_1
Xoutput23 net23 VGND VGND VPWR VPWR prod[15] sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_27_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_643_ _010_ net16 _254_ VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__and3b_1
X_574_ _293_ _007_ _008_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_488_ _236_ _246_ _248_ _249_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__a211o_1
X_626_ net8 VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__inv_2
X_557_ _280_ _304_ _305_ VGND VGND VPWR VPWR _306_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_411_ _143_ _146_ _174_ VGND VGND VPWR VPWR _176_ sky130_fd_sc_hd__nand3_1
X_342_ _094_ _096_ _106_ VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__a21oi_1
X_609_ net51 _042_ _011_ _043_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__o31a_1
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_325_ _088_ _089_ VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_0_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_45 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_590_ _021_ _023_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput24 net24 VGND VGND VPWR VPWR prod[1] sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_642_ net44 net15 VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__nand2_1
X_573_ _297_ _006_ VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_625_ _247_ VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__inv_2
X_487_ _241_ _244_ VGND VGND VPWR VPWR _249_ sky130_fd_sc_hd__or2_1
X_556_ _283_ _286_ VGND VGND VPWR VPWR _305_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_410_ _143_ _146_ _174_ VGND VGND VPWR VPWR _175_ sky130_fd_sc_hd__a21o_1
X_341_ _104_ _105_ VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_0_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_608_ net43 net14 net13 _272_ VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__a22o_1
X_539_ _280_ _287_ VGND VGND VPWR VPWR _288_ sky130_fd_sc_hd__xnor2_1
X_324_ _266_ _265_ VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_13_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_3_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_641_ _040_ _047_ VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__and2b_1
Xoutput25 net25 VGND VGND VPWR VPWR prod[2] sky130_fd_sc_hd__clkbuf_4
X_572_ _297_ _006_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_486_ _228_ _238_ _225_ VGND VGND VPWR VPWR _248_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_555_ _283_ _286_ VGND VGND VPWR VPWR _304_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_624_ _247_ net7 net8 _255_ VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__a22o_1
X_607_ net14 VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__inv_2
X_340_ _100_ _103_ VGND VGND VPWR VPWR _105_ sky130_fd_sc_hd__and2_1
X_538_ _283_ net48 VGND VGND VPWR VPWR _287_ sky130_fd_sc_hd__xnor2_1
X_469_ _214_ _217_ _231_ VGND VGND VPWR VPWR _232_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_13_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_323_ _086_ _087_ VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_112 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_571_ _298_ _005_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__xnor2_1
Xoutput26 net26 VGND VGND VPWR VPWR prod[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_640_ _036_ _073_ _074_ VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__a21o_1
X_485_ _236_ _246_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__xor2_1
XFILLER_0_13_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_554_ _299_ _300_ _302_ VGND VGND VPWR VPWR _303_ sky130_fd_sc_hd__o21ai_1
X_623_ _056_ _057_ VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__or2_1
X_468_ _223_ _230_ VGND VGND VPWR VPWR _231_ sky130_fd_sc_hd__xnor2_1
X_399_ _127_ _129_ _163_ VGND VGND VPWR VPWR _164_ sky130_fd_sc_hd__a21o_1
X_606_ _011_ _294_ _295_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__a21oi_1
X_537_ net47 _285_ VGND VGND VPWR VPWR _286_ sky130_fd_sc_hd__xnor2_1
X_322_ _076_ _049_ _085_ VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__or3_1
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_124 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput27 net27 VGND VGND VPWR VPWR prod[4] sky130_fd_sc_hd__clkbuf_4
X_570_ _303_ _004_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__xor2_1
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_89 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_484_ _244_ _245_ VGND VGND VPWR VPWR _246_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_553_ net35 _301_ _266_ net38 VGND VGND VPWR VPWR _302_ sky130_fd_sc_hd__a22o_1
X_622_ _270_ net6 _023_ VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_19_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_467_ _228_ _229_ VGND VGND VPWR VPWR _230_ sky130_fd_sc_hd__or2_1
X_398_ _161_ _162_ VGND VGND VPWR VPWR _163_ sky130_fd_sc_hd__nand2_1
X_605_ _254_ _037_ _010_ _039_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_536_ _247_ _272_ _258_ VGND VGND VPWR VPWR _285_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_321_ _076_ _049_ _085_ VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_10_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_519_ net2 net12 VGND VGND VPWR VPWR _268_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_7_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput17 net17 VGND VGND VPWR VPWR prod[0] sky130_fd_sc_hd__clkbuf_4
Xoutput28 net28 VGND VGND VPWR VPWR prod[5] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_26_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_483_ _220_ _234_ _243_ VGND VGND VPWR VPWR _245_ sky130_fd_sc_hd__a21oi_1
X_552_ net6 VGND VGND VPWR VPWR _301_ sky130_fd_sc_hd__buf_2
X_621_ _261_ _301_ _266_ _270_ VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_0_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_466_ _224_ _225_ _226_ VGND VGND VPWR VPWR _229_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_397_ _272_ _037_ _123_ VGND VGND VPWR VPWR _162_ sky130_fd_sc_hd__nand3_1
X_604_ _253_ net16 _038_ _254_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__a22oi_1
XPHY_EDGE_ROW_20_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_535_ _273_ _274_ _275_ VGND VGND VPWR VPWR _284_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_320_ _083_ _084_ VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_449_ _101_ net14 _154_ VGND VGND VPWR VPWR _212_ sky130_fd_sc_hd__and3_1
X_518_ net1 _261_ VGND VGND VPWR VPWR _267_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_23_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput18 net18 VGND VGND VPWR VPWR prod[10] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput29 net29 VGND VGND VPWR VPWR prod[6] sky130_fd_sc_hd__buf_2
XFILLER_0_7_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_620_ _030_ _027_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__and2b_1
X_551_ net38 net6 VGND VGND VPWR VPWR _300_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_482_ _220_ _234_ _243_ VGND VGND VPWR VPWR _244_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_20_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_465_ _224_ _225_ _226_ VGND VGND VPWR VPWR _228_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_396_ _272_ _037_ _077_ _123_ VGND VGND VPWR VPWR _161_ sky130_fd_sc_hd__a31o_1
X_603_ net15 VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__buf_2
X_534_ _281_ _282_ VGND VGND VPWR VPWR _283_ sky130_fd_sc_hd__xor2_2
XFILLER_0_4_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_448_ _209_ _210_ VGND VGND VPWR VPWR _211_ sky130_fd_sc_hd__xor2_1
X_379_ _141_ _142_ _137_ VGND VGND VPWR VPWR _144_ sky130_fd_sc_hd__o21ai_1
X_517_ net5 VGND VGND VPWR VPWR _266_ sky130_fd_sc_hd__buf_2
XFILLER_0_5_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput19 net19 VGND VGND VPWR VPWR prod[11] sky130_fd_sc_hd__buf_2
XFILLER_0_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_481_ _241_ _242_ VGND VGND VPWR VPWR _243_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_550_ net34 net5 VGND VGND VPWR VPWR _299_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_20_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_464_ _097_ _038_ _210_ _184_ VGND VGND VPWR VPWR _226_ sky130_fd_sc_hd__a31o_1
X_602_ net16 VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__buf_2
X_533_ _262_ _268_ VGND VGND VPWR VPWR _282_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_395_ _158_ _159_ VGND VGND VPWR VPWR _160_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_447_ _301_ _037_ _157_ VGND VGND VPWR VPWR _210_ sky130_fd_sc_hd__and3_1
X_516_ net13 VGND VGND VPWR VPWR _265_ sky130_fd_sc_hd__buf_2
X_378_ _137_ _141_ _142_ VGND VGND VPWR VPWR _143_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_0_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_480_ _237_ _232_ _240_ VGND VGND VPWR VPWR _242_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_3_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_601_ _009_ _034_ _035_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__a21o_1
X_463_ _097_ _101_ _037_ _038_ VGND VGND VPWR VPWR _225_ sky130_fd_sc_hd__nand4_1
XFILLER_0_24_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_394_ _156_ _157_ VGND VGND VPWR VPWR _159_ sky130_fd_sc_hd__nand2_1
X_532_ net3 net11 VGND VGND VPWR VPWR _281_ sky130_fd_sc_hd__nand2_4
XFILLER_0_14_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_446_ _097_ _038_ VGND VGND VPWR VPWR _209_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_377_ _138_ _139_ _140_ VGND VGND VPWR VPWR _142_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_0_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_515_ _263_ net39 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__nor2_1
XFILLER_0_25_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_104 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_429_ _158_ _192_ VGND VGND VPWR VPWR _193_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput1 a[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_27_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_462_ _097_ _037_ _038_ _101_ VGND VGND VPWR VPWR _224_ sky130_fd_sc_hd__a22o_1
X_393_ _156_ _157_ VGND VGND VPWR VPWR _158_ sky130_fd_sc_hd__or2_1
X_531_ _264_ _278_ _279_ VGND VGND VPWR VPWR _280_ sky130_fd_sc_hd__a21o_1
X_600_ _016_ _033_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_514_ _259_ _260_ _262_ VGND VGND VPWR VPWR _264_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_84 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_445_ _185_ _191_ VGND VGND VPWR VPWR _208_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_376_ _138_ _139_ _140_ VGND VGND VPWR VPWR _141_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_359_ _119_ _121_ _122_ VGND VGND VPWR VPWR _124_ sky130_fd_sc_hd__a21oi_1
X_428_ _185_ _191_ VGND VGND VPWR VPWR _192_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput2 a[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_20_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_461_ _189_ _212_ _187_ VGND VGND VPWR VPWR _223_ sky130_fd_sc_hd__a21bo_1
X_392_ _266_ _038_ VGND VGND VPWR VPWR _157_ sky130_fd_sc_hd__nand2_1
X_530_ _277_ _269_ _271_ _276_ VGND VGND VPWR VPWR _279_ sky130_fd_sc_hd__and4_1
XFILLER_0_14_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_444_ _196_ _195_ VGND VGND VPWR VPWR _207_ sky130_fd_sc_hd__or2b_1
X_375_ _261_ _097_ _099_ _057_ VGND VGND VPWR VPWR _140_ sky130_fd_sc_hd__a31o_1
X_513_ _259_ _260_ _262_ VGND VGND VPWR VPWR _263_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_358_ _119_ _121_ _122_ VGND VGND VPWR VPWR _123_ sky130_fd_sc_hd__and3_1
X_427_ _189_ _190_ VGND VGND VPWR VPWR _191_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 a[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_8
XFILLER_0_11_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_460_ _206_ _222_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__xor2_1
X_391_ _154_ _155_ VGND VGND VPWR VPWR _156_ sky130_fd_sc_hd__xor2_1
XFILLER_0_14_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_589_ _021_ _023_ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__and2_1
X_443_ _181_ _204_ _205_ VGND VGND VPWR VPWR _206_ sky130_fd_sc_hd__a21o_1
X_374_ _309_ _061_ _098_ VGND VGND VPWR VPWR _139_ sky130_fd_sc_hd__or3_1
X_512_ _253_ _261_ VGND VGND VPWR VPWR _262_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_357_ _253_ net45 net16 _038_ _254_ VGND VGND VPWR VPWR _122_ sky130_fd_sc_hd__o2111a_1
X_426_ _186_ _187_ _188_ VGND VGND VPWR VPWR _190_ sky130_fd_sc_hd__a21oi_1
Xinput4 a[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_6
XFILLER_0_22_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_409_ _270_ _101_ _141_ _173_ VGND VGND VPWR VPWR _174_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_124 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_390_ _301_ net14 _089_ VGND VGND VPWR VPWR _155_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_588_ _022_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_18_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_442_ _203_ _200_ VGND VGND VPWR VPWR _205_ sky130_fd_sc_hd__and2b_1
X_373_ _270_ _097_ _101_ _261_ VGND VGND VPWR VPWR _138_ sky130_fd_sc_hd__a22o_1
X_511_ net11 VGND VGND VPWR VPWR _261_ sky130_fd_sc_hd__buf_4
XFILLER_0_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_356_ net52 _120_ _077_ VGND VGND VPWR VPWR _121_ sky130_fd_sc_hd__or3_1
X_425_ _186_ _187_ _188_ VGND VGND VPWR VPWR _189_ sky130_fd_sc_hd__and3_1
Xinput5 a[4] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
XFILLER_0_22_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_408_ _141_ _172_ VGND VGND VPWR VPWR _173_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_339_ _100_ _103_ VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_136 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_6_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_587_ _261_ net5 VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__nand2_1
X_441_ _181_ _204_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__xor2_1
X_372_ _064_ _102_ _062_ VGND VGND VPWR VPWR _137_ sky130_fd_sc_hd__a21boi_1
X_510_ _247_ _254_ _227_ net41 _255_ VGND VGND VPWR VPWR _260_ sky130_fd_sc_hd__a32o_1
X_639_ _051_ _072_ VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_355_ net16 VGND VGND VPWR VPWR _120_ sky130_fd_sc_hd__inv_2
X_424_ _266_ _097_ net14 _265_ _301_ VGND VGND VPWR VPWR _188_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_11_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput6 a[5] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_407_ _270_ _101_ _098_ VGND VGND VPWR VPWR _172_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_338_ _064_ _102_ VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_9 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_586_ _019_ _020_ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__xnor2_1
X_440_ _200_ _203_ VGND VGND VPWR VPWR _204_ sky130_fd_sc_hd__xnor2_1
X_371_ _109_ _093_ VGND VGND VPWR VPWR _136_ sky130_fd_sc_hd__and2b_1
X_569_ _306_ _003_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__xor2_1
X_638_ _051_ _072_ VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_354_ net45 net16 _038_ _272_ VGND VGND VPWR VPWR _119_ sky130_fd_sc_hd__a22o_1
X_423_ _061_ _042_ _154_ VGND VGND VPWR VPWR _187_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_102 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 a[6] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
XFILLER_0_9_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_406_ _136_ _148_ VGND VGND VPWR VPWR _171_ sky130_fd_sc_hd__and2_1
X_337_ _247_ _101_ _019_ VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_25_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput10 b[1] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_4
XFILLER_0_3_146 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_585_ net38 net6 _299_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__and3_1
X_370_ _133_ _134_ VGND VGND VPWR VPWR _135_ sky130_fd_sc_hd__or2_1
X_637_ _053_ _071_ VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__xnor2_2
X_568_ _002_ _001_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__and2_4
XFILLER_0_5_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_499_ _227_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__inv_2
X_422_ _097_ net14 _265_ _101_ VGND VGND VPWR VPWR _186_ sky130_fd_sc_hd__a22o_1
X_353_ net46 _265_ _045_ VGND VGND VPWR VPWR _118_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 a[7] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_1
XFILLER_0_14_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_405_ _168_ _169_ VGND VGND VPWR VPWR _170_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_336_ net8 VGND VGND VPWR VPWR _101_ sky130_fd_sc_hd__buf_2
XFILLER_0_6_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_319_ _079_ _082_ VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__or2_1
Xinput11 b[2] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_4
XFILLER_0_3_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_584_ _255_ net7 VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__nand2_2
XFILLER_0_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_567_ net33 _000_ _307_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__o21ai_1
X_636_ _069_ _070_ VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__or2b_4
X_498_ net1 net9 VGND VGND VPWR VPWR _227_ sky130_fd_sc_hd__nand2_1
X_421_ _183_ _184_ VGND VGND VPWR VPWR _185_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_14_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_352_ _114_ _116_ VGND VGND VPWR VPWR _117_ sky130_fd_sc_hd__nand2_1
Xinput9 b[0] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
X_619_ _257_ _261_ _272_ _270_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_404_ _153_ _133_ _167_ VGND VGND VPWR VPWR _169_ sky130_fd_sc_hd__nor3_1
X_335_ _098_ _099_ VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_318_ _079_ _082_ VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput12 b[3] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_10_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_80 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_583_ _298_ _005_ _017_ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_9 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_497_ net40 _252_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__xnor2_1
X_566_ _307_ _313_ _000_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__or3_4
X_635_ _068_ _054_ _028_ _055_ VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_14_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_420_ _301_ _266_ _037_ _038_ VGND VGND VPWR VPWR _184_ sky130_fd_sc_hd__and4_1
X_351_ _115_ _042_ _089_ VGND VGND VPWR VPWR _116_ sky130_fd_sc_hd__or3_1
XFILLER_0_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_549_ _289_ VGND VGND VPWR VPWR _298_ sky130_fd_sc_hd__inv_2
X_618_ _018_ _032_ _052_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_403_ _153_ _133_ _167_ VGND VGND VPWR VPWR _168_ sky130_fd_sc_hd__o21a_1
X_334_ _270_ _301_ _022_ VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_317_ _045_ _081_ VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__xor2_1
Xinput13 b[4] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
XFILLER_0_23_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_582_ _303_ _004_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__or2b_1
XFILLER_0_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_496_ _279_ _278_ VGND VGND VPWR VPWR _252_ sky130_fd_sc_hd__or2b_1
X_634_ _054_ _028_ _055_ _068_ VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__o31a_1
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_565_ _310_ _311_ _312_ VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_350_ _301_ VGND VGND VPWR VPWR _115_ sky130_fd_sc_hd__inv_2
X_479_ _237_ _232_ _240_ VGND VGND VPWR VPWR _241_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_548_ _294_ _295_ _296_ VGND VGND VPWR VPWR _297_ sky130_fd_sc_hd__o21ai_2
X_617_ _026_ _031_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_402_ _160_ _166_ VGND VGND VPWR VPWR _167_ sky130_fd_sc_hd__xor2_1
X_333_ _261_ _097_ VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput14 b[5] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_2
X_316_ _011_ _080_ VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_581_ _014_ _015_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_495_ _292_ _250_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__nor2_1
X_564_ _310_ _311_ _312_ VGND VGND VPWR VPWR _313_ sky130_fd_sc_hd__and3_1
X_633_ _024_ _067_ VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_83 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_478_ _101_ _037_ _228_ _239_ VGND VGND VPWR VPWR _240_ sky130_fd_sc_hd__a31o_1
X_616_ _049_ _050_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__nor2_1
X_547_ _253_ net14 _265_ _254_ VGND VGND VPWR VPWR _296_ sky130_fd_sc_hd__a22o_1
X_401_ _164_ _165_ VGND VGND VPWR VPWR _166_ sky130_fd_sc_hd__nand2_1
X_332_ net7 VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_11_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput15 b[6] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_1
X_315_ net52 _042_ VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_580_ _010_ _013_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_563_ _267_ _281_ _268_ VGND VGND VPWR VPWR _312_ sky130_fd_sc_hd__a21oi_1
X_632_ _058_ _066_ VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_95 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_494_ _253_ _265_ _291_ VGND VGND VPWR VPWR _250_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_477_ _228_ _238_ VGND VGND VPWR VPWR _239_ sky130_fd_sc_hd__nor2_1
X_615_ _014_ _048_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__and2_1
X_546_ _254_ net14 VGND VGND VPWR VPWR _295_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_400_ _127_ _129_ _163_ VGND VGND VPWR VPWR _165_ sky130_fd_sc_hd__nand3_1
XFILLER_0_6_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_331_ _024_ _095_ VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_529_ _269_ _271_ _276_ _277_ VGND VGND VPWR VPWR _278_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput16 b[7] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
X_314_ _077_ _078_ VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__xor2_1
XFILLER_0_23_40 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_493_ _113_ _150_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__xor2_1
X_562_ _261_ _272_ net12 _257_ VGND VGND VPWR VPWR _311_ sky130_fd_sc_hd__a22o_1
X_631_ _064_ _065_ VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_476_ _101_ _037_ _209_ VGND VGND VPWR VPWR _238_ sky130_fd_sc_hd__and3_1
X_614_ _014_ _048_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__nor2_1
X_545_ _253_ _265_ VGND VGND VPWR VPWR _294_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_330_ _067_ VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__inv_2
X_459_ _220_ _221_ VGND VGND VPWR VPWR _222_ sky130_fd_sc_hd__nor2_1
X_528_ _273_ _274_ _275_ VGND VGND VPWR VPWR _277_ sky130_fd_sc_hd__nand3_1
XFILLER_0_10_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_561_ _308_ _309_ _281_ VGND VGND VPWR VPWR _310_ sky130_fd_sc_hd__or3_4
X_630_ _059_ _062_ _063_ VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__a21oi_1
X_492_ _075_ _111_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__xor2_1
XFILLER_0_17_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_613_ _040_ _047_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__xor2_1
X_475_ _230_ _223_ VGND VGND VPWR VPWR _237_ sky130_fd_sc_hd__or2b_1
XFILLER_0_26_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_544_ _292_ VGND VGND VPWR VPWR _293_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_458_ _207_ _198_ _219_ VGND VGND VPWR VPWR _221_ sky130_fd_sc_hd__and3_1
X_389_ _097_ _265_ VGND VGND VPWR VPWR _154_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_527_ _273_ _274_ _275_ VGND VGND VPWR VPWR _276_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_21_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_491_ _036_ _073_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__xor2_1
X_560_ net12 VGND VGND VPWR VPWR _309_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_474_ _206_ _222_ _234_ VGND VGND VPWR VPWR _236_ sky130_fd_sc_hd__and3_1
X_612_ _045_ _046_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__nor2_1
X_543_ _253_ _265_ _291_ VGND VGND VPWR VPWR _292_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_526_ net1 net3 net2 net10 net9 VGND VGND VPWR VPWR _275_ sky130_fd_sc_hd__o2111a_1
X_457_ _207_ _198_ _219_ VGND VGND VPWR VPWR _220_ sky130_fd_sc_hd__a21oi_2
X_388_ _114_ _116_ _131_ VGND VGND VPWR VPWR _153_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_509_ _251_ _258_ _227_ VGND VGND VPWR VPWR _259_ sky130_fd_sc_hd__or3b_4
XTAP_TAPCELL_ROW_21_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_490_ _009_ _034_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__xor2_1
XFILLER_0_9_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_473_ _234_ _235_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__xnor2_1
X_611_ _041_ _044_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__nor2_1
X_542_ _289_ _290_ VGND VGND VPWR VPWR _291_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer20 net51 VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_8_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_456_ _217_ _218_ VGND VGND VPWR VPWR _219_ sky130_fd_sc_hd__or2_1
X_387_ _113_ _150_ _151_ VGND VGND VPWR VPWR _152_ sky130_fd_sc_hd__a21o_1
X_525_ net10 net3 net4 net9 VGND VGND VPWR VPWR _274_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_439_ _175_ _201_ _202_ VGND VGND VPWR VPWR _203_ sky130_fd_sc_hd__and3_1
X_508_ _255_ _257_ VGND VGND VPWR VPWR _258_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_25_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_44 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_472_ _206_ _222_ _220_ VGND VGND VPWR VPWR _235_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_610_ _041_ _044_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__and2_1
X_541_ net37 _266_ _288_ VGND VGND VPWR VPWR _290_ sky130_fd_sc_hd__a21oi_1
Xrebuffer10 _257_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_27_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_455_ _208_ _193_ _216_ VGND VGND VPWR VPWR _218_ sky130_fd_sc_hd__and3_1
X_386_ _135_ _149_ VGND VGND VPWR VPWR _151_ sky130_fd_sc_hd__nor2_1
X_524_ _255_ net10 net3 _272_ VGND VGND VPWR VPWR _273_ sky130_fd_sc_hd__nand4_2
XFILLER_0_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_369_ _090_ _132_ VGND VGND VPWR VPWR _134_ sky130_fd_sc_hd__and2_1
X_438_ _141_ _172_ _139_ VGND VGND VPWR VPWR _202_ sky130_fd_sc_hd__a21boi_1
Xrebuffer1 net50 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
X_507_ net3 VGND VGND VPWR VPWR _257_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_5_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_471_ _232_ _233_ VGND VGND VPWR VPWR _234_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_540_ net36 _266_ _288_ VGND VGND VPWR VPWR _289_ sky130_fd_sc_hd__and3_1
Xrebuffer11 net42 VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_454_ _208_ _193_ _216_ VGND VGND VPWR VPWR _217_ sky130_fd_sc_hd__a21oi_1
X_385_ _135_ _149_ VGND VGND VPWR VPWR _150_ sky130_fd_sc_hd__xor2_1
X_523_ net4 VGND VGND VPWR VPWR _272_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_368_ _090_ _132_ VGND VGND VPWR VPWR _133_ sky130_fd_sc_hd__nor2_1
X_437_ _171_ _177_ VGND VGND VPWR VPWR _201_ sky130_fd_sc_hd__nand2_1
Xrebuffer2 _255_ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
X_506_ _227_ _251_ _256_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__o21a_1
XFILLER_0_18_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_470_ _214_ _217_ _231_ VGND VGND VPWR VPWR _233_ sky130_fd_sc_hd__or3_1
X_599_ _016_ _033_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__xor2_1
Xrebuffer12 net42 VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_1
XFILLER_0_13_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_453_ _214_ _215_ VGND VGND VPWR VPWR _216_ sky130_fd_sc_hd__or2_1
X_384_ _136_ _148_ VGND VGND VPWR VPWR _149_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_12_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_522_ _254_ _261_ _270_ _253_ VGND VGND VPWR VPWR _271_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_436_ _198_ _199_ VGND VGND VPWR VPWR _200_ sky130_fd_sc_hd__and2_1
X_367_ _117_ _131_ VGND VGND VPWR VPWR _132_ sky130_fd_sc_hd__xor2_1
XFILLER_0_2_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer3 net34 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_1
X_505_ _253_ _247_ _254_ _255_ VGND VGND VPWR VPWR _256_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_58 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_419_ _266_ _037_ _038_ _301_ VGND VGND VPWR VPWR _183_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer13 net44 VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_16_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_598_ _018_ _032_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__xor2_1
X_452_ _211_ _213_ VGND VGND VPWR VPWR _215_ sky130_fd_sc_hd__and2_1
X_383_ _146_ _147_ VGND VGND VPWR VPWR _148_ sky130_fd_sc_hd__and2_1
X_521_ net12 VGND VGND VPWR VPWR _270_ sky130_fd_sc_hd__buf_2
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_435_ _182_ _168_ _197_ VGND VGND VPWR VPWR _199_ sky130_fd_sc_hd__or3_1
X_366_ _129_ _130_ VGND VGND VPWR VPWR _131_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer4 net35 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
X_504_ net9 VGND VGND VPWR VPWR _255_ sky130_fd_sc_hd__buf_6
XFILLER_0_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_418_ _160_ _166_ VGND VGND VPWR VPWR _182_ sky130_fd_sc_hd__nor2_1
X_349_ _266_ net14 _265_ _301_ VGND VGND VPWR VPWR _114_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_597_ _026_ _031_ VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer14 net44 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_520_ _267_ _268_ VGND VGND VPWR VPWR _269_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_451_ _211_ _213_ VGND VGND VPWR VPWR _214_ sky130_fd_sc_hd__nor2_1
X_382_ _104_ _107_ _145_ VGND VGND VPWR VPWR _147_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_2_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_136 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_434_ _182_ _168_ _197_ VGND VGND VPWR VPWR _198_ sky130_fd_sc_hd__o21ai_2
X_365_ _084_ _086_ _128_ VGND VGND VPWR VPWR _130_ sky130_fd_sc_hd__nand3_1
X_503_ net2 VGND VGND VPWR VPWR _254_ sky130_fd_sc_hd__buf_2
XFILLER_0_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer5 net36 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_417_ _152_ _179_ _180_ VGND VGND VPWR VPWR _181_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_348_ _075_ _111_ _112_ VGND VGND VPWR VPWR _113_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_596_ net49 _030_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_15_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer15 _284_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_450_ _189_ _212_ VGND VGND VPWR VPWR _213_ sky130_fd_sc_hd__xnor2_1
X_381_ _104_ _107_ _145_ VGND VGND VPWR VPWR _146_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_579_ _010_ _013_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_433_ _195_ _196_ VGND VGND VPWR VPWR _197_ sky130_fd_sc_hd__xnor2_1
X_502_ net1 VGND VGND VPWR VPWR _253_ sky130_fd_sc_hd__buf_2
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_364_ _084_ _086_ _128_ VGND VGND VPWR VPWR _129_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer6 _247_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_1
X_416_ _170_ _178_ VGND VGND VPWR VPWR _180_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_347_ _092_ _110_ VGND VGND VPWR VPWR _112_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_595_ _028_ _029_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__or2b_1
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer16 _286_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_380_ _143_ _144_ VGND VGND VPWR VPWR _145_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput30 net30 VGND VGND VPWR VPWR prod[7] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_18_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_578_ _011_ _012_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__xnor2_1
.ends

